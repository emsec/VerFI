
module Cipher ( clk, rst, Input, Key, Output, done );
  input [63:0] Input;
  input [127:0] Key;
  output [63:0] Output;
  input clk, rst;
  output done;
  wire   RoundConstant_4_, RoundConstant_0, selects_0_, selectsReg_0_,
         selectsNext_0_, MCInst_XOR_r0_Inst_0_n5, MCInst_XOR_r0_Inst_1_n5,
         MCInst_XOR_r0_Inst_2_n5, MCInst_XOR_r0_Inst_3_n5,
         MCInst_XOR_r0_Inst_4_n5, MCInst_XOR_r0_Inst_5_n5,
         MCInst_XOR_r0_Inst_6_n5, MCInst_XOR_r0_Inst_7_n5,
         MCInst_XOR_r0_Inst_8_n5, MCInst_XOR_r0_Inst_9_n5,
         MCInst_XOR_r0_Inst_10_n5, MCInst_XOR_r0_Inst_11_n5,
         MCInst_XOR_r0_Inst_12_n5, MCInst_XOR_r0_Inst_13_n5,
         MCInst_XOR_r0_Inst_14_n5, MCInst_XOR_r0_Inst_15_n5,
         AddKeyConstXOR_XORInst_0_0_n5, AddKeyConstXOR_XORInst_0_1_n5,
         AddKeyConstXOR_XORInst_0_2_n5, AddKeyConstXOR_XORInst_1_0_n5,
         AddKeyConstXOR_XORInst_1_1_n5, AddKeyConstXOR_XORInst_1_2_n5,
         AddKeyConstXOR_XORInst_1_3_n5, SubCellInst_LFInst_0_n7,
         SubCellInst_LFInst_0_n6, SubCellInst_LFInst_0_n5,
         SubCellInst_LFInst_0_n4, SubCellInst_LFInst_0_n3,
         SubCellInst_LFInst_0_n2, SubCellInst_LFInst_0_n1,
         SubCellInst_LFInst_1_n27, SubCellInst_LFInst_1_n26,
         SubCellInst_LFInst_1_n25, SubCellInst_LFInst_1_n24,
         SubCellInst_LFInst_1_n23, SubCellInst_LFInst_1_n22,
         SubCellInst_LFInst_1_n21, SubCellInst_LFInst_2_n27,
         SubCellInst_LFInst_2_n26, SubCellInst_LFInst_2_n25,
         SubCellInst_LFInst_2_n24, SubCellInst_LFInst_2_n23,
         SubCellInst_LFInst_2_n22, SubCellInst_LFInst_2_n21,
         SubCellInst_LFInst_3_n27, SubCellInst_LFInst_3_n26,
         SubCellInst_LFInst_3_n25, SubCellInst_LFInst_3_n24,
         SubCellInst_LFInst_3_n23, SubCellInst_LFInst_3_n22,
         SubCellInst_LFInst_3_n21, SubCellInst_LFInst_4_n27,
         SubCellInst_LFInst_4_n26, SubCellInst_LFInst_4_n25,
         SubCellInst_LFInst_4_n24, SubCellInst_LFInst_4_n23,
         SubCellInst_LFInst_4_n22, SubCellInst_LFInst_4_n21,
         SubCellInst_LFInst_5_n27, SubCellInst_LFInst_5_n26,
         SubCellInst_LFInst_5_n25, SubCellInst_LFInst_5_n24,
         SubCellInst_LFInst_5_n23, SubCellInst_LFInst_5_n22,
         SubCellInst_LFInst_5_n21, SubCellInst_LFInst_6_n27,
         SubCellInst_LFInst_6_n26, SubCellInst_LFInst_6_n25,
         SubCellInst_LFInst_6_n24, SubCellInst_LFInst_6_n23,
         SubCellInst_LFInst_6_n22, SubCellInst_LFInst_6_n21,
         SubCellInst_LFInst_7_n27, SubCellInst_LFInst_7_n26,
         SubCellInst_LFInst_7_n25, SubCellInst_LFInst_7_n24,
         SubCellInst_LFInst_7_n23, SubCellInst_LFInst_7_n22,
         SubCellInst_LFInst_7_n21, SubCellInst_LFInst_8_n27,
         SubCellInst_LFInst_8_n26, SubCellInst_LFInst_8_n25,
         SubCellInst_LFInst_8_n24, SubCellInst_LFInst_8_n23,
         SubCellInst_LFInst_8_n22, SubCellInst_LFInst_8_n21,
         SubCellInst_LFInst_9_n27, SubCellInst_LFInst_9_n26,
         SubCellInst_LFInst_9_n25, SubCellInst_LFInst_9_n24,
         SubCellInst_LFInst_9_n23, SubCellInst_LFInst_9_n22,
         SubCellInst_LFInst_9_n21, SubCellInst_LFInst_10_n27,
         SubCellInst_LFInst_10_n26, SubCellInst_LFInst_10_n25,
         SubCellInst_LFInst_10_n24, SubCellInst_LFInst_10_n23,
         SubCellInst_LFInst_10_n22, SubCellInst_LFInst_10_n21,
         SubCellInst_LFInst_11_n27, SubCellInst_LFInst_11_n26,
         SubCellInst_LFInst_11_n25, SubCellInst_LFInst_11_n24,
         SubCellInst_LFInst_11_n23, SubCellInst_LFInst_11_n22,
         SubCellInst_LFInst_11_n21, SubCellInst_LFInst_12_n27,
         SubCellInst_LFInst_12_n26, SubCellInst_LFInst_12_n25,
         SubCellInst_LFInst_12_n24, SubCellInst_LFInst_12_n23,
         SubCellInst_LFInst_12_n22, SubCellInst_LFInst_12_n21,
         SubCellInst_LFInst_13_n27, SubCellInst_LFInst_13_n26,
         SubCellInst_LFInst_13_n25, SubCellInst_LFInst_13_n24,
         SubCellInst_LFInst_13_n23, SubCellInst_LFInst_13_n22,
         SubCellInst_LFInst_13_n21, SubCellInst_LFInst_14_n27,
         SubCellInst_LFInst_14_n26, SubCellInst_LFInst_14_n25,
         SubCellInst_LFInst_14_n24, SubCellInst_LFInst_14_n23,
         SubCellInst_LFInst_14_n22, SubCellInst_LFInst_14_n21,
         SubCellInst_LFInst_15_n27, SubCellInst_LFInst_15_n26,
         SubCellInst_LFInst_15_n25, SubCellInst_LFInst_15_n24,
         SubCellInst_LFInst_15_n23, SubCellInst_LFInst_15_n22,
         SubCellInst_LFInst_15_n21, KeyMUX_n7, KeyMUX_n6, KeyMUX_n5,
         FSMMUX_MUXInst_1_n4, FSMMUX_MUXInst_2_n4, FSMMUX_MUXInst_4_n4,
         FSMMUX_MUXInst_5_n4, FSMMUX_MUXInst_6_n4, FSMSignalsInst_n1;
  wire   [63:0] Feedback;
  wire   [63:32] MCInput;
  wire   [63:0] MCOutput;
  wire   [63:0] AddRoundKeyOutput;
  wire   [63:0] SelectedKey;
  wire   [6:0] FSMReg;
  wire   [6:0] FSMUpdate;

  MUX2_X1 InputMUX_MUXInst_0_U1 ( .A(Feedback[0]), .B(Input[0]), .S(rst), .Z(
        MCOutput[0]) );
  MUX2_X1 InputMUX_MUXInst_1_U1 ( .A(Feedback[1]), .B(Input[1]), .S(rst), .Z(
        MCOutput[1]) );
  MUX2_X1 InputMUX_MUXInst_2_U1 ( .A(Feedback[2]), .B(Input[2]), .S(rst), .Z(
        MCOutput[2]) );
  MUX2_X1 InputMUX_MUXInst_3_U1 ( .A(Feedback[3]), .B(Input[3]), .S(rst), .Z(
        MCOutput[3]) );
  MUX2_X1 InputMUX_MUXInst_4_U1 ( .A(Feedback[4]), .B(Input[4]), .S(rst), .Z(
        MCOutput[4]) );
  MUX2_X1 InputMUX_MUXInst_5_U1 ( .A(Feedback[5]), .B(Input[5]), .S(rst), .Z(
        MCOutput[5]) );
  MUX2_X1 InputMUX_MUXInst_6_U1 ( .A(Feedback[6]), .B(Input[6]), .S(rst), .Z(
        MCOutput[6]) );
  MUX2_X1 InputMUX_MUXInst_7_U1 ( .A(Feedback[7]), .B(Input[7]), .S(rst), .Z(
        MCOutput[7]) );
  MUX2_X1 InputMUX_MUXInst_8_U1 ( .A(Feedback[8]), .B(Input[8]), .S(rst), .Z(
        MCOutput[8]) );
  MUX2_X1 InputMUX_MUXInst_9_U1 ( .A(Feedback[9]), .B(Input[9]), .S(rst), .Z(
        MCOutput[9]) );
  MUX2_X1 InputMUX_MUXInst_10_U1 ( .A(Feedback[10]), .B(Input[10]), .S(rst), 
        .Z(MCOutput[10]) );
  MUX2_X1 InputMUX_MUXInst_11_U1 ( .A(Feedback[11]), .B(Input[11]), .S(rst), 
        .Z(MCOutput[11]) );
  MUX2_X1 InputMUX_MUXInst_12_U1 ( .A(Feedback[12]), .B(Input[12]), .S(rst), 
        .Z(MCOutput[12]) );
  MUX2_X1 InputMUX_MUXInst_13_U1 ( .A(Feedback[13]), .B(Input[13]), .S(rst), 
        .Z(MCOutput[13]) );
  MUX2_X1 InputMUX_MUXInst_14_U1 ( .A(Feedback[14]), .B(Input[14]), .S(rst), 
        .Z(MCOutput[14]) );
  MUX2_X1 InputMUX_MUXInst_15_U1 ( .A(Feedback[15]), .B(Input[15]), .S(rst), 
        .Z(MCOutput[15]) );
  MUX2_X1 InputMUX_MUXInst_16_U1 ( .A(Feedback[16]), .B(Input[16]), .S(rst), 
        .Z(MCOutput[16]) );
  MUX2_X1 InputMUX_MUXInst_17_U1 ( .A(Feedback[17]), .B(Input[17]), .S(rst), 
        .Z(MCOutput[17]) );
  MUX2_X1 InputMUX_MUXInst_18_U1 ( .A(Feedback[18]), .B(Input[18]), .S(rst), 
        .Z(MCOutput[18]) );
  MUX2_X1 InputMUX_MUXInst_19_U1 ( .A(Feedback[19]), .B(Input[19]), .S(rst), 
        .Z(MCOutput[19]) );
  MUX2_X1 InputMUX_MUXInst_20_U1 ( .A(Feedback[20]), .B(Input[20]), .S(rst), 
        .Z(MCOutput[20]) );
  MUX2_X1 InputMUX_MUXInst_21_U1 ( .A(Feedback[21]), .B(Input[21]), .S(rst), 
        .Z(MCOutput[21]) );
  MUX2_X1 InputMUX_MUXInst_22_U1 ( .A(Feedback[22]), .B(Input[22]), .S(rst), 
        .Z(MCOutput[22]) );
  MUX2_X1 InputMUX_MUXInst_23_U1 ( .A(Feedback[23]), .B(Input[23]), .S(rst), 
        .Z(MCOutput[23]) );
  MUX2_X1 InputMUX_MUXInst_24_U1 ( .A(Feedback[24]), .B(Input[24]), .S(rst), 
        .Z(MCOutput[24]) );
  MUX2_X1 InputMUX_MUXInst_25_U1 ( .A(Feedback[25]), .B(Input[25]), .S(rst), 
        .Z(MCOutput[25]) );
  MUX2_X1 InputMUX_MUXInst_26_U1 ( .A(Feedback[26]), .B(Input[26]), .S(rst), 
        .Z(MCOutput[26]) );
  MUX2_X1 InputMUX_MUXInst_27_U1 ( .A(Feedback[27]), .B(Input[27]), .S(rst), 
        .Z(MCOutput[27]) );
  MUX2_X1 InputMUX_MUXInst_28_U1 ( .A(Feedback[28]), .B(Input[28]), .S(rst), 
        .Z(MCOutput[28]) );
  MUX2_X1 InputMUX_MUXInst_29_U1 ( .A(Feedback[29]), .B(Input[29]), .S(rst), 
        .Z(MCOutput[29]) );
  MUX2_X1 InputMUX_MUXInst_30_U1 ( .A(Feedback[30]), .B(Input[30]), .S(rst), 
        .Z(MCOutput[30]) );
  MUX2_X1 InputMUX_MUXInst_31_U1 ( .A(Feedback[31]), .B(Input[31]), .S(rst), 
        .Z(MCOutput[31]) );
  MUX2_X1 InputMUX_MUXInst_32_U1 ( .A(Feedback[32]), .B(Input[32]), .S(rst), 
        .Z(MCInput[32]) );
  MUX2_X1 InputMUX_MUXInst_33_U1 ( .A(Feedback[33]), .B(Input[33]), .S(rst), 
        .Z(MCInput[33]) );
  MUX2_X1 InputMUX_MUXInst_34_U1 ( .A(Feedback[34]), .B(Input[34]), .S(rst), 
        .Z(MCInput[34]) );
  MUX2_X1 InputMUX_MUXInst_35_U1 ( .A(Feedback[35]), .B(Input[35]), .S(rst), 
        .Z(MCInput[35]) );
  MUX2_X1 InputMUX_MUXInst_36_U1 ( .A(Feedback[36]), .B(Input[36]), .S(rst), 
        .Z(MCInput[36]) );
  MUX2_X1 InputMUX_MUXInst_37_U1 ( .A(Feedback[37]), .B(Input[37]), .S(rst), 
        .Z(MCInput[37]) );
  MUX2_X1 InputMUX_MUXInst_38_U1 ( .A(Feedback[38]), .B(Input[38]), .S(rst), 
        .Z(MCInput[38]) );
  MUX2_X1 InputMUX_MUXInst_39_U1 ( .A(Feedback[39]), .B(Input[39]), .S(rst), 
        .Z(MCInput[39]) );
  MUX2_X1 InputMUX_MUXInst_40_U1 ( .A(Feedback[40]), .B(Input[40]), .S(rst), 
        .Z(MCInput[40]) );
  MUX2_X1 InputMUX_MUXInst_41_U1 ( .A(Feedback[41]), .B(Input[41]), .S(rst), 
        .Z(MCInput[41]) );
  MUX2_X1 InputMUX_MUXInst_42_U1 ( .A(Feedback[42]), .B(Input[42]), .S(rst), 
        .Z(MCInput[42]) );
  MUX2_X1 InputMUX_MUXInst_43_U1 ( .A(Feedback[43]), .B(Input[43]), .S(rst), 
        .Z(MCInput[43]) );
  MUX2_X1 InputMUX_MUXInst_44_U1 ( .A(Feedback[44]), .B(Input[44]), .S(rst), 
        .Z(MCInput[44]) );
  MUX2_X1 InputMUX_MUXInst_45_U1 ( .A(Feedback[45]), .B(Input[45]), .S(rst), 
        .Z(MCInput[45]) );
  MUX2_X1 InputMUX_MUXInst_46_U1 ( .A(Feedback[46]), .B(Input[46]), .S(rst), 
        .Z(MCInput[46]) );
  MUX2_X1 InputMUX_MUXInst_47_U1 ( .A(Feedback[47]), .B(Input[47]), .S(rst), 
        .Z(MCInput[47]) );
  MUX2_X1 InputMUX_MUXInst_48_U1 ( .A(Feedback[48]), .B(Input[48]), .S(rst), 
        .Z(MCInput[48]) );
  MUX2_X1 InputMUX_MUXInst_49_U1 ( .A(Feedback[49]), .B(Input[49]), .S(rst), 
        .Z(MCInput[49]) );
  MUX2_X1 InputMUX_MUXInst_50_U1 ( .A(Feedback[50]), .B(Input[50]), .S(rst), 
        .Z(MCInput[50]) );
  MUX2_X1 InputMUX_MUXInst_51_U1 ( .A(Feedback[51]), .B(Input[51]), .S(rst), 
        .Z(MCInput[51]) );
  MUX2_X1 InputMUX_MUXInst_52_U1 ( .A(Feedback[52]), .B(Input[52]), .S(rst), 
        .Z(MCInput[52]) );
  MUX2_X1 InputMUX_MUXInst_53_U1 ( .A(Feedback[53]), .B(Input[53]), .S(rst), 
        .Z(MCInput[53]) );
  MUX2_X1 InputMUX_MUXInst_54_U1 ( .A(Feedback[54]), .B(Input[54]), .S(rst), 
        .Z(MCInput[54]) );
  MUX2_X1 InputMUX_MUXInst_55_U1 ( .A(Feedback[55]), .B(Input[55]), .S(rst), 
        .Z(MCInput[55]) );
  MUX2_X1 InputMUX_MUXInst_56_U1 ( .A(Feedback[56]), .B(Input[56]), .S(rst), 
        .Z(MCInput[56]) );
  MUX2_X1 InputMUX_MUXInst_57_U1 ( .A(Feedback[57]), .B(Input[57]), .S(rst), 
        .Z(MCInput[57]) );
  MUX2_X1 InputMUX_MUXInst_58_U1 ( .A(Feedback[58]), .B(Input[58]), .S(rst), 
        .Z(MCInput[58]) );
  MUX2_X1 InputMUX_MUXInst_59_U1 ( .A(Feedback[59]), .B(Input[59]), .S(rst), 
        .Z(MCInput[59]) );
  MUX2_X1 InputMUX_MUXInst_60_U1 ( .A(Feedback[60]), .B(Input[60]), .S(rst), 
        .Z(MCInput[60]) );
  MUX2_X1 InputMUX_MUXInst_61_U1 ( .A(Feedback[61]), .B(Input[61]), .S(rst), 
        .Z(MCInput[61]) );
  MUX2_X1 InputMUX_MUXInst_62_U1 ( .A(Feedback[62]), .B(Input[62]), .S(rst), 
        .Z(MCInput[62]) );
  MUX2_X1 InputMUX_MUXInst_63_U1 ( .A(Feedback[63]), .B(Input[63]), .S(rst), 
        .Z(MCInput[63]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_0_U2 ( .A(MCInst_XOR_r0_Inst_0_n5), .B(
        MCOutput[16]), .ZN(MCOutput[48]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_0_U1 ( .A(MCOutput[0]), .B(MCInput[48]), .ZN(
        MCInst_XOR_r0_Inst_0_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_0_U1 ( .A(MCInput[32]), .B(MCOutput[0]), .Z(
        MCOutput[32]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U2 ( .A(MCInst_XOR_r0_Inst_1_n5), .B(
        MCOutput[17]), .ZN(MCOutput[49]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U1 ( .A(MCOutput[1]), .B(MCInput[49]), .ZN(
        MCInst_XOR_r0_Inst_1_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_1_U1 ( .A(MCInput[33]), .B(MCOutput[1]), .Z(
        MCOutput[33]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U2 ( .A(MCInst_XOR_r0_Inst_2_n5), .B(
        MCOutput[18]), .ZN(MCOutput[50]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U1 ( .A(MCOutput[2]), .B(MCInput[50]), .ZN(
        MCInst_XOR_r0_Inst_2_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_2_U1 ( .A(MCInput[34]), .B(MCOutput[2]), .Z(
        MCOutput[34]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U2 ( .A(MCInst_XOR_r0_Inst_3_n5), .B(
        MCOutput[19]), .ZN(MCOutput[51]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U1 ( .A(MCOutput[3]), .B(MCInput[51]), .ZN(
        MCInst_XOR_r0_Inst_3_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_3_U1 ( .A(MCInput[35]), .B(MCOutput[3]), .Z(
        MCOutput[35]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U2 ( .A(MCInst_XOR_r0_Inst_4_n5), .B(
        MCOutput[20]), .ZN(MCOutput[52]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U1 ( .A(MCOutput[4]), .B(MCInput[52]), .ZN(
        MCInst_XOR_r0_Inst_4_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_4_U1 ( .A(MCInput[36]), .B(MCOutput[4]), .Z(
        MCOutput[36]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U2 ( .A(MCInst_XOR_r0_Inst_5_n5), .B(
        MCOutput[21]), .ZN(MCOutput[53]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U1 ( .A(MCOutput[5]), .B(MCInput[53]), .ZN(
        MCInst_XOR_r0_Inst_5_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_5_U1 ( .A(MCInput[37]), .B(MCOutput[5]), .Z(
        MCOutput[37]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U2 ( .A(MCInst_XOR_r0_Inst_6_n5), .B(
        MCOutput[22]), .ZN(MCOutput[54]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U1 ( .A(MCOutput[6]), .B(MCInput[54]), .ZN(
        MCInst_XOR_r0_Inst_6_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_6_U1 ( .A(MCInput[38]), .B(MCOutput[6]), .Z(
        MCOutput[38]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U2 ( .A(MCInst_XOR_r0_Inst_7_n5), .B(
        MCOutput[23]), .ZN(MCOutput[55]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U1 ( .A(MCOutput[7]), .B(MCInput[55]), .ZN(
        MCInst_XOR_r0_Inst_7_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_7_U1 ( .A(MCInput[39]), .B(MCOutput[7]), .Z(
        MCOutput[39]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U2 ( .A(MCInst_XOR_r0_Inst_8_n5), .B(
        MCOutput[24]), .ZN(MCOutput[56]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U1 ( .A(MCOutput[8]), .B(MCInput[56]), .ZN(
        MCInst_XOR_r0_Inst_8_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_8_U1 ( .A(MCInput[40]), .B(MCOutput[8]), .Z(
        MCOutput[40]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U2 ( .A(MCInst_XOR_r0_Inst_9_n5), .B(
        MCOutput[25]), .ZN(MCOutput[57]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U1 ( .A(MCOutput[9]), .B(MCInput[57]), .ZN(
        MCInst_XOR_r0_Inst_9_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_9_U1 ( .A(MCInput[41]), .B(MCOutput[9]), .Z(
        MCOutput[41]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U2 ( .A(MCInst_XOR_r0_Inst_10_n5), .B(
        MCOutput[26]), .ZN(MCOutput[58]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U1 ( .A(MCOutput[10]), .B(MCInput[58]), .ZN(
        MCInst_XOR_r0_Inst_10_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_10_U1 ( .A(MCInput[42]), .B(MCOutput[10]), .Z(
        MCOutput[42]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U2 ( .A(MCInst_XOR_r0_Inst_11_n5), .B(
        MCOutput[27]), .ZN(MCOutput[59]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U1 ( .A(MCOutput[11]), .B(MCInput[59]), .ZN(
        MCInst_XOR_r0_Inst_11_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_11_U1 ( .A(MCInput[43]), .B(MCOutput[11]), .Z(
        MCOutput[43]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U2 ( .A(MCInst_XOR_r0_Inst_12_n5), .B(
        MCOutput[28]), .ZN(MCOutput[60]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U1 ( .A(MCOutput[12]), .B(MCInput[60]), .ZN(
        MCInst_XOR_r0_Inst_12_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_12_U1 ( .A(MCInput[44]), .B(MCOutput[12]), .Z(
        MCOutput[44]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U2 ( .A(MCInst_XOR_r0_Inst_13_n5), .B(
        MCOutput[29]), .ZN(MCOutput[61]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U1 ( .A(MCOutput[13]), .B(MCInput[61]), .ZN(
        MCInst_XOR_r0_Inst_13_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_13_U1 ( .A(MCInput[45]), .B(MCOutput[13]), .Z(
        MCOutput[45]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U2 ( .A(MCInst_XOR_r0_Inst_14_n5), .B(
        MCOutput[30]), .ZN(MCOutput[62]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U1 ( .A(MCOutput[14]), .B(MCInput[62]), .ZN(
        MCInst_XOR_r0_Inst_14_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_14_U1 ( .A(MCInput[46]), .B(MCOutput[14]), .Z(
        MCOutput[46]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U2 ( .A(MCInst_XOR_r0_Inst_15_n5), .B(
        MCOutput[31]), .ZN(MCOutput[63]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U1 ( .A(MCOutput[15]), .B(MCInput[63]), .ZN(
        MCInst_XOR_r0_Inst_15_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_15_U1 ( .A(MCInput[47]), .B(MCOutput[15]), .Z(
        MCOutput[47]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_0_U1 ( .A(MCOutput[48]), .B(SelectedKey[48]), 
        .Z(AddRoundKeyOutput[48]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_1_U1 ( .A(MCOutput[49]), .B(SelectedKey[49]), 
        .Z(AddRoundKeyOutput[49]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_2_U1 ( .A(MCOutput[50]), .B(SelectedKey[50]), 
        .Z(AddRoundKeyOutput[50]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_3_U1 ( .A(MCOutput[51]), .B(SelectedKey[51]), 
        .Z(AddRoundKeyOutput[51]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_0_U1 ( .A(MCOutput[52]), .B(SelectedKey[52]), 
        .Z(AddRoundKeyOutput[52]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_1_U1 ( .A(MCOutput[53]), .B(SelectedKey[53]), 
        .Z(AddRoundKeyOutput[53]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_2_U1 ( .A(MCOutput[54]), .B(SelectedKey[54]), 
        .Z(AddRoundKeyOutput[54]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_3_U1 ( .A(MCOutput[55]), .B(SelectedKey[55]), 
        .Z(AddRoundKeyOutput[55]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_0_U1 ( .A(MCOutput[56]), .B(SelectedKey[56]), 
        .Z(AddRoundKeyOutput[56]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_1_U1 ( .A(MCOutput[57]), .B(SelectedKey[57]), 
        .Z(AddRoundKeyOutput[57]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_2_U1 ( .A(MCOutput[58]), .B(SelectedKey[58]), 
        .Z(AddRoundKeyOutput[58]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_3_U1 ( .A(MCOutput[59]), .B(SelectedKey[59]), 
        .Z(AddRoundKeyOutput[59]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_0_U1 ( .A(MCOutput[60]), .B(SelectedKey[60]), 
        .Z(AddRoundKeyOutput[60]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_1_U1 ( .A(MCOutput[61]), .B(SelectedKey[61]), 
        .Z(AddRoundKeyOutput[61]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_2_U1 ( .A(MCOutput[62]), .B(SelectedKey[62]), 
        .Z(AddRoundKeyOutput[62]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_3_U1 ( .A(MCOutput[63]), .B(SelectedKey[63]), 
        .Z(AddRoundKeyOutput[63]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_0_U2 ( .A(AddKeyConstXOR_XORInst_0_0_n5), 
        .B(SelectedKey[40]), .ZN(AddRoundKeyOutput[40]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_0_U1 ( .A(RoundConstant_0), .B(
        MCOutput[40]), .ZN(AddKeyConstXOR_XORInst_0_0_n5) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_1_U2 ( .A(AddKeyConstXOR_XORInst_0_1_n5), 
        .B(SelectedKey[41]), .ZN(AddRoundKeyOutput[41]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_1_U1 ( .A(FSMUpdate[0]), .B(MCOutput[41]), 
        .ZN(AddKeyConstXOR_XORInst_0_1_n5) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_2_U2 ( .A(AddKeyConstXOR_XORInst_0_2_n5), 
        .B(SelectedKey[42]), .ZN(AddRoundKeyOutput[42]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_2_U1 ( .A(FSMUpdate[1]), .B(MCOutput[42]), 
        .ZN(AddKeyConstXOR_XORInst_0_2_n5) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_3_U1 ( .A(MCOutput[43]), .B(SelectedKey[43]), .Z(AddRoundKeyOutput[43]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_0_U2 ( .A(AddKeyConstXOR_XORInst_1_0_n5), 
        .B(SelectedKey[44]), .ZN(AddRoundKeyOutput[44]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_0_U1 ( .A(RoundConstant_4_), .B(
        MCOutput[44]), .ZN(AddKeyConstXOR_XORInst_1_0_n5) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_1_U2 ( .A(AddKeyConstXOR_XORInst_1_1_n5), 
        .B(SelectedKey[45]), .ZN(AddRoundKeyOutput[45]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_1_U1 ( .A(FSMUpdate[3]), .B(MCOutput[45]), 
        .ZN(AddKeyConstXOR_XORInst_1_1_n5) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_2_U2 ( .A(AddKeyConstXOR_XORInst_1_2_n5), 
        .B(SelectedKey[46]), .ZN(AddRoundKeyOutput[46]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_2_U1 ( .A(FSMUpdate[4]), .B(MCOutput[46]), 
        .ZN(AddKeyConstXOR_XORInst_1_2_n5) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_3_U2 ( .A(AddKeyConstXOR_XORInst_1_3_n5), 
        .B(SelectedKey[47]), .ZN(AddRoundKeyOutput[47]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_3_U1 ( .A(FSMUpdate[5]), .B(MCOutput[47]), 
        .ZN(AddKeyConstXOR_XORInst_1_3_n5) );
  XOR2_X1 AddKeyXOR2_XORInst_0_0_U1 ( .A(MCOutput[0]), .B(SelectedKey[0]), .Z(
        AddRoundKeyOutput[0]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_1_U1 ( .A(MCOutput[1]), .B(SelectedKey[1]), .Z(
        AddRoundKeyOutput[1]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_2_U1 ( .A(MCOutput[2]), .B(SelectedKey[2]), .Z(
        AddRoundKeyOutput[2]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_3_U1 ( .A(MCOutput[3]), .B(SelectedKey[3]), .Z(
        AddRoundKeyOutput[3]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_0_U1 ( .A(MCOutput[4]), .B(SelectedKey[4]), .Z(
        AddRoundKeyOutput[4]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_1_U1 ( .A(MCOutput[5]), .B(SelectedKey[5]), .Z(
        AddRoundKeyOutput[5]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_2_U1 ( .A(MCOutput[6]), .B(SelectedKey[6]), .Z(
        AddRoundKeyOutput[6]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_3_U1 ( .A(MCOutput[7]), .B(SelectedKey[7]), .Z(
        AddRoundKeyOutput[7]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_0_U1 ( .A(MCOutput[8]), .B(SelectedKey[8]), .Z(
        AddRoundKeyOutput[8]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_1_U1 ( .A(MCOutput[9]), .B(SelectedKey[9]), .Z(
        AddRoundKeyOutput[9]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_2_U1 ( .A(MCOutput[10]), .B(SelectedKey[10]), 
        .Z(AddRoundKeyOutput[10]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_3_U1 ( .A(MCOutput[11]), .B(SelectedKey[11]), 
        .Z(AddRoundKeyOutput[11]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_0_U1 ( .A(MCOutput[12]), .B(SelectedKey[12]), 
        .Z(AddRoundKeyOutput[12]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_1_U1 ( .A(MCOutput[13]), .B(SelectedKey[13]), 
        .Z(AddRoundKeyOutput[13]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_2_U1 ( .A(MCOutput[14]), .B(SelectedKey[14]), 
        .Z(AddRoundKeyOutput[14]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_3_U1 ( .A(MCOutput[15]), .B(SelectedKey[15]), 
        .Z(AddRoundKeyOutput[15]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_0_U1 ( .A(MCOutput[16]), .B(SelectedKey[16]), 
        .Z(AddRoundKeyOutput[16]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_1_U1 ( .A(MCOutput[17]), .B(SelectedKey[17]), 
        .Z(AddRoundKeyOutput[17]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_2_U1 ( .A(MCOutput[18]), .B(SelectedKey[18]), 
        .Z(AddRoundKeyOutput[18]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_3_U1 ( .A(MCOutput[19]), .B(SelectedKey[19]), 
        .Z(AddRoundKeyOutput[19]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_0_U1 ( .A(MCOutput[20]), .B(SelectedKey[20]), 
        .Z(AddRoundKeyOutput[20]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_1_U1 ( .A(MCOutput[21]), .B(SelectedKey[21]), 
        .Z(AddRoundKeyOutput[21]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_2_U1 ( .A(MCOutput[22]), .B(SelectedKey[22]), 
        .Z(AddRoundKeyOutput[22]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_3_U1 ( .A(MCOutput[23]), .B(SelectedKey[23]), 
        .Z(AddRoundKeyOutput[23]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_0_U1 ( .A(MCOutput[24]), .B(SelectedKey[24]), 
        .Z(AddRoundKeyOutput[24]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_1_U1 ( .A(MCOutput[25]), .B(SelectedKey[25]), 
        .Z(AddRoundKeyOutput[25]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_2_U1 ( .A(MCOutput[26]), .B(SelectedKey[26]), 
        .Z(AddRoundKeyOutput[26]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_3_U1 ( .A(MCOutput[27]), .B(SelectedKey[27]), 
        .Z(AddRoundKeyOutput[27]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_0_U1 ( .A(MCOutput[28]), .B(SelectedKey[28]), 
        .Z(AddRoundKeyOutput[28]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_1_U1 ( .A(MCOutput[29]), .B(SelectedKey[29]), 
        .Z(AddRoundKeyOutput[29]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_2_U1 ( .A(MCOutput[30]), .B(SelectedKey[30]), 
        .Z(AddRoundKeyOutput[30]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_3_U1 ( .A(MCOutput[31]), .B(SelectedKey[31]), 
        .Z(AddRoundKeyOutput[31]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_0_U1 ( .A(MCOutput[32]), .B(SelectedKey[32]), 
        .Z(AddRoundKeyOutput[32]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_1_U1 ( .A(MCOutput[33]), .B(SelectedKey[33]), 
        .Z(AddRoundKeyOutput[33]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_2_U1 ( .A(MCOutput[34]), .B(SelectedKey[34]), 
        .Z(AddRoundKeyOutput[34]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_3_U1 ( .A(MCOutput[35]), .B(SelectedKey[35]), 
        .Z(AddRoundKeyOutput[35]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_0_U1 ( .A(MCOutput[36]), .B(SelectedKey[36]), 
        .Z(AddRoundKeyOutput[36]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_1_U1 ( .A(MCOutput[37]), .B(SelectedKey[37]), 
        .Z(AddRoundKeyOutput[37]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_2_U1 ( .A(MCOutput[38]), .B(SelectedKey[38]), 
        .Z(AddRoundKeyOutput[38]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_3_U1 ( .A(MCOutput[39]), .B(SelectedKey[39]), 
        .Z(AddRoundKeyOutput[39]) );
  DFF_X1 StateReg_s_current_state_reg_0_ ( .D(AddRoundKeyOutput[0]), .CK(clk), 
        .Q(Output[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1_ ( .D(AddRoundKeyOutput[1]), .CK(clk), 
        .Q(Output[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2_ ( .D(AddRoundKeyOutput[2]), .CK(clk), 
        .Q(Output[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3_ ( .D(AddRoundKeyOutput[3]), .CK(clk), 
        .Q(Output[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4_ ( .D(AddRoundKeyOutput[4]), .CK(clk), 
        .Q(Output[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5_ ( .D(AddRoundKeyOutput[5]), .CK(clk), 
        .Q(Output[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6_ ( .D(AddRoundKeyOutput[6]), .CK(clk), 
        .Q(Output[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7_ ( .D(AddRoundKeyOutput[7]), .CK(clk), 
        .Q(Output[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8_ ( .D(AddRoundKeyOutput[8]), .CK(clk), 
        .Q(Output[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9_ ( .D(AddRoundKeyOutput[9]), .CK(clk), 
        .Q(Output[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10_ ( .D(AddRoundKeyOutput[10]), .CK(clk), .Q(Output[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11_ ( .D(AddRoundKeyOutput[11]), .CK(clk), .Q(Output[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12_ ( .D(AddRoundKeyOutput[12]), .CK(clk), .Q(Output[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13_ ( .D(AddRoundKeyOutput[13]), .CK(clk), .Q(Output[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14_ ( .D(AddRoundKeyOutput[14]), .CK(clk), .Q(Output[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15_ ( .D(AddRoundKeyOutput[15]), .CK(clk), .Q(Output[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16_ ( .D(AddRoundKeyOutput[16]), .CK(clk), .Q(Output[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17_ ( .D(AddRoundKeyOutput[17]), .CK(clk), .Q(Output[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18_ ( .D(AddRoundKeyOutput[18]), .CK(clk), .Q(Output[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19_ ( .D(AddRoundKeyOutput[19]), .CK(clk), .Q(Output[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20_ ( .D(AddRoundKeyOutput[20]), .CK(clk), .Q(Output[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21_ ( .D(AddRoundKeyOutput[21]), .CK(clk), .Q(Output[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22_ ( .D(AddRoundKeyOutput[22]), .CK(clk), .Q(Output[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23_ ( .D(AddRoundKeyOutput[23]), .CK(clk), .Q(Output[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24_ ( .D(AddRoundKeyOutput[24]), .CK(clk), .Q(Output[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25_ ( .D(AddRoundKeyOutput[25]), .CK(clk), .Q(Output[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26_ ( .D(AddRoundKeyOutput[26]), .CK(clk), .Q(Output[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27_ ( .D(AddRoundKeyOutput[27]), .CK(clk), .Q(Output[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28_ ( .D(AddRoundKeyOutput[28]), .CK(clk), .Q(Output[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29_ ( .D(AddRoundKeyOutput[29]), .CK(clk), .Q(Output[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30_ ( .D(AddRoundKeyOutput[30]), .CK(clk), .Q(Output[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31_ ( .D(AddRoundKeyOutput[31]), .CK(clk), .Q(Output[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32_ ( .D(AddRoundKeyOutput[32]), .CK(clk), .Q(Output[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33_ ( .D(AddRoundKeyOutput[33]), .CK(clk), .Q(Output[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34_ ( .D(AddRoundKeyOutput[34]), .CK(clk), .Q(Output[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35_ ( .D(AddRoundKeyOutput[35]), .CK(clk), .Q(Output[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36_ ( .D(AddRoundKeyOutput[36]), .CK(clk), .Q(Output[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37_ ( .D(AddRoundKeyOutput[37]), .CK(clk), .Q(Output[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38_ ( .D(AddRoundKeyOutput[38]), .CK(clk), .Q(Output[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39_ ( .D(AddRoundKeyOutput[39]), .CK(clk), .Q(Output[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40_ ( .D(AddRoundKeyOutput[40]), .CK(clk), .Q(Output[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41_ ( .D(AddRoundKeyOutput[41]), .CK(clk), .Q(Output[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42_ ( .D(AddRoundKeyOutput[42]), .CK(clk), .Q(Output[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43_ ( .D(AddRoundKeyOutput[43]), .CK(clk), .Q(Output[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44_ ( .D(AddRoundKeyOutput[44]), .CK(clk), .Q(Output[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45_ ( .D(AddRoundKeyOutput[45]), .CK(clk), .Q(Output[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46_ ( .D(AddRoundKeyOutput[46]), .CK(clk), .Q(Output[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47_ ( .D(AddRoundKeyOutput[47]), .CK(clk), .Q(Output[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48_ ( .D(AddRoundKeyOutput[48]), .CK(clk), .Q(Output[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49_ ( .D(AddRoundKeyOutput[49]), .CK(clk), .Q(Output[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50_ ( .D(AddRoundKeyOutput[50]), .CK(clk), .Q(Output[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51_ ( .D(AddRoundKeyOutput[51]), .CK(clk), .Q(Output[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52_ ( .D(AddRoundKeyOutput[52]), .CK(clk), .Q(Output[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53_ ( .D(AddRoundKeyOutput[53]), .CK(clk), .Q(Output[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54_ ( .D(AddRoundKeyOutput[54]), .CK(clk), .Q(Output[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55_ ( .D(AddRoundKeyOutput[55]), .CK(clk), .Q(Output[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56_ ( .D(AddRoundKeyOutput[56]), .CK(clk), .Q(Output[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57_ ( .D(AddRoundKeyOutput[57]), .CK(clk), .Q(Output[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58_ ( .D(AddRoundKeyOutput[58]), .CK(clk), .Q(Output[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59_ ( .D(AddRoundKeyOutput[59]), .CK(clk), .Q(Output[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60_ ( .D(AddRoundKeyOutput[60]), .CK(clk), .Q(Output[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61_ ( .D(AddRoundKeyOutput[61]), .CK(clk), .Q(Output[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62_ ( .D(AddRoundKeyOutput[62]), .CK(clk), .Q(Output[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63_ ( .D(AddRoundKeyOutput[63]), .CK(clk), .Q(Output[63]), .QN() );
  OAI22_X1 SubCellInst_LFInst_0_U11 ( .A1(Output[63]), .A2(Output[60]), .B1(
        SubCellInst_LFInst_0_n7), .B2(Output[61]), .ZN(Feedback[3]) );
  NOR2_X1 SubCellInst_LFInst_0_U10 ( .A1(SubCellInst_LFInst_0_n6), .A2(
        SubCellInst_LFInst_0_n5), .ZN(SubCellInst_LFInst_0_n7) );
  OAI22_X1 SubCellInst_LFInst_0_U9 ( .A1(Output[63]), .A2(Output[60]), .B1(
        SubCellInst_LFInst_0_n4), .B2(SubCellInst_LFInst_0_n3), .ZN(
        Feedback[2]) );
  AOI21_X1 SubCellInst_LFInst_0_U8 ( .B1(Output[60]), .B2(Output[63]), .A(
        Output[62]), .ZN(SubCellInst_LFInst_0_n3) );
  OAI21_X1 SubCellInst_LFInst_0_U7 ( .B1(Output[63]), .B2(
        SubCellInst_LFInst_0_n6), .A(SubCellInst_LFInst_0_n2), .ZN(Feedback[1]) );
  OAI21_X1 SubCellInst_LFInst_0_U6 ( .B1(Output[62]), .B2(
        SubCellInst_LFInst_0_n5), .A(Output[60]), .ZN(SubCellInst_LFInst_0_n2)
         );
  INV_X1 SubCellInst_LFInst_0_U5 ( .A(Output[63]), .ZN(SubCellInst_LFInst_0_n5) );
  INV_X1 SubCellInst_LFInst_0_U4 ( .A(Output[62]), .ZN(SubCellInst_LFInst_0_n6) );
  AOI22_X1 SubCellInst_LFInst_0_U3 ( .A1(Output[63]), .A2(Output[62]), .B1(
        SubCellInst_LFInst_0_n1), .B2(SubCellInst_LFInst_0_n4), .ZN(
        Feedback[0]) );
  INV_X1 SubCellInst_LFInst_0_U2 ( .A(Output[61]), .ZN(SubCellInst_LFInst_0_n4) );
  OAI21_X1 SubCellInst_LFInst_0_U1 ( .B1(Output[62]), .B2(Output[63]), .A(
        Output[60]), .ZN(SubCellInst_LFInst_0_n1) );
  OAI22_X1 SubCellInst_LFInst_1_U11 ( .A1(Output[51]), .A2(Output[48]), .B1(
        SubCellInst_LFInst_1_n27), .B2(Output[49]), .ZN(Feedback[7]) );
  NOR2_X1 SubCellInst_LFInst_1_U10 ( .A1(SubCellInst_LFInst_1_n26), .A2(
        SubCellInst_LFInst_1_n25), .ZN(SubCellInst_LFInst_1_n27) );
  OAI22_X1 SubCellInst_LFInst_1_U9 ( .A1(Output[51]), .A2(Output[48]), .B1(
        SubCellInst_LFInst_1_n24), .B2(SubCellInst_LFInst_1_n23), .ZN(
        Feedback[6]) );
  AOI21_X1 SubCellInst_LFInst_1_U8 ( .B1(Output[48]), .B2(Output[51]), .A(
        Output[50]), .ZN(SubCellInst_LFInst_1_n23) );
  OAI21_X1 SubCellInst_LFInst_1_U7 ( .B1(Output[51]), .B2(
        SubCellInst_LFInst_1_n26), .A(SubCellInst_LFInst_1_n22), .ZN(
        Feedback[5]) );
  OAI21_X1 SubCellInst_LFInst_1_U6 ( .B1(Output[50]), .B2(
        SubCellInst_LFInst_1_n25), .A(Output[48]), .ZN(
        SubCellInst_LFInst_1_n22) );
  INV_X1 SubCellInst_LFInst_1_U5 ( .A(Output[51]), .ZN(
        SubCellInst_LFInst_1_n25) );
  INV_X1 SubCellInst_LFInst_1_U4 ( .A(Output[50]), .ZN(
        SubCellInst_LFInst_1_n26) );
  AOI22_X1 SubCellInst_LFInst_1_U3 ( .A1(Output[51]), .A2(Output[50]), .B1(
        SubCellInst_LFInst_1_n21), .B2(SubCellInst_LFInst_1_n24), .ZN(
        Feedback[4]) );
  INV_X1 SubCellInst_LFInst_1_U2 ( .A(Output[49]), .ZN(
        SubCellInst_LFInst_1_n24) );
  OAI21_X1 SubCellInst_LFInst_1_U1 ( .B1(Output[50]), .B2(Output[51]), .A(
        Output[48]), .ZN(SubCellInst_LFInst_1_n21) );
  OAI22_X1 SubCellInst_LFInst_2_U11 ( .A1(Output[55]), .A2(Output[52]), .B1(
        SubCellInst_LFInst_2_n27), .B2(Output[53]), .ZN(Feedback[11]) );
  NOR2_X1 SubCellInst_LFInst_2_U10 ( .A1(SubCellInst_LFInst_2_n26), .A2(
        SubCellInst_LFInst_2_n25), .ZN(SubCellInst_LFInst_2_n27) );
  OAI22_X1 SubCellInst_LFInst_2_U9 ( .A1(Output[55]), .A2(Output[52]), .B1(
        SubCellInst_LFInst_2_n24), .B2(SubCellInst_LFInst_2_n23), .ZN(
        Feedback[10]) );
  AOI21_X1 SubCellInst_LFInst_2_U8 ( .B1(Output[52]), .B2(Output[55]), .A(
        Output[54]), .ZN(SubCellInst_LFInst_2_n23) );
  OAI21_X1 SubCellInst_LFInst_2_U7 ( .B1(Output[55]), .B2(
        SubCellInst_LFInst_2_n26), .A(SubCellInst_LFInst_2_n22), .ZN(
        Feedback[9]) );
  OAI21_X1 SubCellInst_LFInst_2_U6 ( .B1(Output[54]), .B2(
        SubCellInst_LFInst_2_n25), .A(Output[52]), .ZN(
        SubCellInst_LFInst_2_n22) );
  INV_X1 SubCellInst_LFInst_2_U5 ( .A(Output[55]), .ZN(
        SubCellInst_LFInst_2_n25) );
  INV_X1 SubCellInst_LFInst_2_U4 ( .A(Output[54]), .ZN(
        SubCellInst_LFInst_2_n26) );
  AOI22_X1 SubCellInst_LFInst_2_U3 ( .A1(Output[55]), .A2(Output[54]), .B1(
        SubCellInst_LFInst_2_n21), .B2(SubCellInst_LFInst_2_n24), .ZN(
        Feedback[8]) );
  INV_X1 SubCellInst_LFInst_2_U2 ( .A(Output[53]), .ZN(
        SubCellInst_LFInst_2_n24) );
  OAI21_X1 SubCellInst_LFInst_2_U1 ( .B1(Output[54]), .B2(Output[55]), .A(
        Output[52]), .ZN(SubCellInst_LFInst_2_n21) );
  OAI22_X1 SubCellInst_LFInst_3_U11 ( .A1(Output[59]), .A2(Output[56]), .B1(
        SubCellInst_LFInst_3_n27), .B2(Output[57]), .ZN(Feedback[15]) );
  NOR2_X1 SubCellInst_LFInst_3_U10 ( .A1(SubCellInst_LFInst_3_n26), .A2(
        SubCellInst_LFInst_3_n25), .ZN(SubCellInst_LFInst_3_n27) );
  OAI22_X1 SubCellInst_LFInst_3_U9 ( .A1(Output[59]), .A2(Output[56]), .B1(
        SubCellInst_LFInst_3_n24), .B2(SubCellInst_LFInst_3_n23), .ZN(
        Feedback[14]) );
  AOI21_X1 SubCellInst_LFInst_3_U8 ( .B1(Output[56]), .B2(Output[59]), .A(
        Output[58]), .ZN(SubCellInst_LFInst_3_n23) );
  OAI21_X1 SubCellInst_LFInst_3_U7 ( .B1(Output[59]), .B2(
        SubCellInst_LFInst_3_n26), .A(SubCellInst_LFInst_3_n22), .ZN(
        Feedback[13]) );
  OAI21_X1 SubCellInst_LFInst_3_U6 ( .B1(Output[58]), .B2(
        SubCellInst_LFInst_3_n25), .A(Output[56]), .ZN(
        SubCellInst_LFInst_3_n22) );
  INV_X1 SubCellInst_LFInst_3_U5 ( .A(Output[59]), .ZN(
        SubCellInst_LFInst_3_n25) );
  INV_X1 SubCellInst_LFInst_3_U4 ( .A(Output[58]), .ZN(
        SubCellInst_LFInst_3_n26) );
  AOI22_X1 SubCellInst_LFInst_3_U3 ( .A1(Output[59]), .A2(Output[58]), .B1(
        SubCellInst_LFInst_3_n21), .B2(SubCellInst_LFInst_3_n24), .ZN(
        Feedback[12]) );
  INV_X1 SubCellInst_LFInst_3_U2 ( .A(Output[57]), .ZN(
        SubCellInst_LFInst_3_n24) );
  OAI21_X1 SubCellInst_LFInst_3_U1 ( .B1(Output[58]), .B2(Output[59]), .A(
        Output[56]), .ZN(SubCellInst_LFInst_3_n21) );
  OAI22_X1 SubCellInst_LFInst_4_U11 ( .A1(Output[35]), .A2(Output[32]), .B1(
        SubCellInst_LFInst_4_n27), .B2(Output[33]), .ZN(Feedback[19]) );
  NOR2_X1 SubCellInst_LFInst_4_U10 ( .A1(SubCellInst_LFInst_4_n26), .A2(
        SubCellInst_LFInst_4_n25), .ZN(SubCellInst_LFInst_4_n27) );
  OAI22_X1 SubCellInst_LFInst_4_U9 ( .A1(Output[35]), .A2(Output[32]), .B1(
        SubCellInst_LFInst_4_n24), .B2(SubCellInst_LFInst_4_n23), .ZN(
        Feedback[18]) );
  AOI21_X1 SubCellInst_LFInst_4_U8 ( .B1(Output[32]), .B2(Output[35]), .A(
        Output[34]), .ZN(SubCellInst_LFInst_4_n23) );
  OAI21_X1 SubCellInst_LFInst_4_U7 ( .B1(Output[35]), .B2(
        SubCellInst_LFInst_4_n26), .A(SubCellInst_LFInst_4_n22), .ZN(
        Feedback[17]) );
  OAI21_X1 SubCellInst_LFInst_4_U6 ( .B1(Output[34]), .B2(
        SubCellInst_LFInst_4_n25), .A(Output[32]), .ZN(
        SubCellInst_LFInst_4_n22) );
  INV_X1 SubCellInst_LFInst_4_U5 ( .A(Output[35]), .ZN(
        SubCellInst_LFInst_4_n25) );
  INV_X1 SubCellInst_LFInst_4_U4 ( .A(Output[34]), .ZN(
        SubCellInst_LFInst_4_n26) );
  AOI22_X1 SubCellInst_LFInst_4_U3 ( .A1(Output[35]), .A2(Output[34]), .B1(
        SubCellInst_LFInst_4_n21), .B2(SubCellInst_LFInst_4_n24), .ZN(
        Feedback[16]) );
  INV_X1 SubCellInst_LFInst_4_U2 ( .A(Output[33]), .ZN(
        SubCellInst_LFInst_4_n24) );
  OAI21_X1 SubCellInst_LFInst_4_U1 ( .B1(Output[34]), .B2(Output[35]), .A(
        Output[32]), .ZN(SubCellInst_LFInst_4_n21) );
  OAI22_X1 SubCellInst_LFInst_5_U11 ( .A1(Output[47]), .A2(Output[44]), .B1(
        SubCellInst_LFInst_5_n27), .B2(Output[45]), .ZN(Feedback[23]) );
  NOR2_X1 SubCellInst_LFInst_5_U10 ( .A1(SubCellInst_LFInst_5_n26), .A2(
        SubCellInst_LFInst_5_n25), .ZN(SubCellInst_LFInst_5_n27) );
  OAI22_X1 SubCellInst_LFInst_5_U9 ( .A1(Output[47]), .A2(Output[44]), .B1(
        SubCellInst_LFInst_5_n24), .B2(SubCellInst_LFInst_5_n23), .ZN(
        Feedback[22]) );
  AOI21_X1 SubCellInst_LFInst_5_U8 ( .B1(Output[44]), .B2(Output[47]), .A(
        Output[46]), .ZN(SubCellInst_LFInst_5_n23) );
  OAI21_X1 SubCellInst_LFInst_5_U7 ( .B1(Output[47]), .B2(
        SubCellInst_LFInst_5_n26), .A(SubCellInst_LFInst_5_n22), .ZN(
        Feedback[21]) );
  OAI21_X1 SubCellInst_LFInst_5_U6 ( .B1(Output[46]), .B2(
        SubCellInst_LFInst_5_n25), .A(Output[44]), .ZN(
        SubCellInst_LFInst_5_n22) );
  INV_X1 SubCellInst_LFInst_5_U5 ( .A(Output[47]), .ZN(
        SubCellInst_LFInst_5_n25) );
  INV_X1 SubCellInst_LFInst_5_U4 ( .A(Output[46]), .ZN(
        SubCellInst_LFInst_5_n26) );
  AOI22_X1 SubCellInst_LFInst_5_U3 ( .A1(Output[47]), .A2(Output[46]), .B1(
        SubCellInst_LFInst_5_n21), .B2(SubCellInst_LFInst_5_n24), .ZN(
        Feedback[20]) );
  INV_X1 SubCellInst_LFInst_5_U2 ( .A(Output[45]), .ZN(
        SubCellInst_LFInst_5_n24) );
  OAI21_X1 SubCellInst_LFInst_5_U1 ( .B1(Output[46]), .B2(Output[47]), .A(
        Output[44]), .ZN(SubCellInst_LFInst_5_n21) );
  OAI22_X1 SubCellInst_LFInst_6_U11 ( .A1(Output[43]), .A2(Output[40]), .B1(
        SubCellInst_LFInst_6_n27), .B2(Output[41]), .ZN(Feedback[27]) );
  NOR2_X1 SubCellInst_LFInst_6_U10 ( .A1(SubCellInst_LFInst_6_n26), .A2(
        SubCellInst_LFInst_6_n25), .ZN(SubCellInst_LFInst_6_n27) );
  OAI22_X1 SubCellInst_LFInst_6_U9 ( .A1(Output[43]), .A2(Output[40]), .B1(
        SubCellInst_LFInst_6_n24), .B2(SubCellInst_LFInst_6_n23), .ZN(
        Feedback[26]) );
  AOI21_X1 SubCellInst_LFInst_6_U8 ( .B1(Output[40]), .B2(Output[43]), .A(
        Output[42]), .ZN(SubCellInst_LFInst_6_n23) );
  OAI21_X1 SubCellInst_LFInst_6_U7 ( .B1(Output[43]), .B2(
        SubCellInst_LFInst_6_n26), .A(SubCellInst_LFInst_6_n22), .ZN(
        Feedback[25]) );
  OAI21_X1 SubCellInst_LFInst_6_U6 ( .B1(Output[42]), .B2(
        SubCellInst_LFInst_6_n25), .A(Output[40]), .ZN(
        SubCellInst_LFInst_6_n22) );
  INV_X1 SubCellInst_LFInst_6_U5 ( .A(Output[43]), .ZN(
        SubCellInst_LFInst_6_n25) );
  INV_X1 SubCellInst_LFInst_6_U4 ( .A(Output[42]), .ZN(
        SubCellInst_LFInst_6_n26) );
  AOI22_X1 SubCellInst_LFInst_6_U3 ( .A1(Output[43]), .A2(Output[42]), .B1(
        SubCellInst_LFInst_6_n21), .B2(SubCellInst_LFInst_6_n24), .ZN(
        Feedback[24]) );
  INV_X1 SubCellInst_LFInst_6_U2 ( .A(Output[41]), .ZN(
        SubCellInst_LFInst_6_n24) );
  OAI21_X1 SubCellInst_LFInst_6_U1 ( .B1(Output[42]), .B2(Output[43]), .A(
        Output[40]), .ZN(SubCellInst_LFInst_6_n21) );
  OAI22_X1 SubCellInst_LFInst_7_U11 ( .A1(Output[39]), .A2(Output[36]), .B1(
        SubCellInst_LFInst_7_n27), .B2(Output[37]), .ZN(Feedback[31]) );
  NOR2_X1 SubCellInst_LFInst_7_U10 ( .A1(SubCellInst_LFInst_7_n26), .A2(
        SubCellInst_LFInst_7_n25), .ZN(SubCellInst_LFInst_7_n27) );
  OAI22_X1 SubCellInst_LFInst_7_U9 ( .A1(Output[39]), .A2(Output[36]), .B1(
        SubCellInst_LFInst_7_n24), .B2(SubCellInst_LFInst_7_n23), .ZN(
        Feedback[30]) );
  AOI21_X1 SubCellInst_LFInst_7_U8 ( .B1(Output[36]), .B2(Output[39]), .A(
        Output[38]), .ZN(SubCellInst_LFInst_7_n23) );
  OAI21_X1 SubCellInst_LFInst_7_U7 ( .B1(Output[39]), .B2(
        SubCellInst_LFInst_7_n26), .A(SubCellInst_LFInst_7_n22), .ZN(
        Feedback[29]) );
  OAI21_X1 SubCellInst_LFInst_7_U6 ( .B1(Output[38]), .B2(
        SubCellInst_LFInst_7_n25), .A(Output[36]), .ZN(
        SubCellInst_LFInst_7_n22) );
  INV_X1 SubCellInst_LFInst_7_U5 ( .A(Output[39]), .ZN(
        SubCellInst_LFInst_7_n25) );
  INV_X1 SubCellInst_LFInst_7_U4 ( .A(Output[38]), .ZN(
        SubCellInst_LFInst_7_n26) );
  AOI22_X1 SubCellInst_LFInst_7_U3 ( .A1(Output[39]), .A2(Output[38]), .B1(
        SubCellInst_LFInst_7_n21), .B2(SubCellInst_LFInst_7_n24), .ZN(
        Feedback[28]) );
  INV_X1 SubCellInst_LFInst_7_U2 ( .A(Output[37]), .ZN(
        SubCellInst_LFInst_7_n24) );
  OAI21_X1 SubCellInst_LFInst_7_U1 ( .B1(Output[38]), .B2(Output[39]), .A(
        Output[36]), .ZN(SubCellInst_LFInst_7_n21) );
  OAI22_X1 SubCellInst_LFInst_8_U11 ( .A1(Output[19]), .A2(Output[16]), .B1(
        SubCellInst_LFInst_8_n27), .B2(Output[17]), .ZN(Feedback[35]) );
  NOR2_X1 SubCellInst_LFInst_8_U10 ( .A1(SubCellInst_LFInst_8_n26), .A2(
        SubCellInst_LFInst_8_n25), .ZN(SubCellInst_LFInst_8_n27) );
  OAI22_X1 SubCellInst_LFInst_8_U9 ( .A1(Output[19]), .A2(Output[16]), .B1(
        SubCellInst_LFInst_8_n24), .B2(SubCellInst_LFInst_8_n23), .ZN(
        Feedback[34]) );
  AOI21_X1 SubCellInst_LFInst_8_U8 ( .B1(Output[16]), .B2(Output[19]), .A(
        Output[18]), .ZN(SubCellInst_LFInst_8_n23) );
  OAI21_X1 SubCellInst_LFInst_8_U7 ( .B1(Output[19]), .B2(
        SubCellInst_LFInst_8_n26), .A(SubCellInst_LFInst_8_n22), .ZN(
        Feedback[33]) );
  OAI21_X1 SubCellInst_LFInst_8_U6 ( .B1(Output[18]), .B2(
        SubCellInst_LFInst_8_n25), .A(Output[16]), .ZN(
        SubCellInst_LFInst_8_n22) );
  INV_X1 SubCellInst_LFInst_8_U5 ( .A(Output[19]), .ZN(
        SubCellInst_LFInst_8_n25) );
  INV_X1 SubCellInst_LFInst_8_U4 ( .A(Output[18]), .ZN(
        SubCellInst_LFInst_8_n26) );
  AOI22_X1 SubCellInst_LFInst_8_U3 ( .A1(Output[19]), .A2(Output[18]), .B1(
        SubCellInst_LFInst_8_n21), .B2(SubCellInst_LFInst_8_n24), .ZN(
        Feedback[32]) );
  INV_X1 SubCellInst_LFInst_8_U2 ( .A(Output[17]), .ZN(
        SubCellInst_LFInst_8_n24) );
  OAI21_X1 SubCellInst_LFInst_8_U1 ( .B1(Output[18]), .B2(Output[19]), .A(
        Output[16]), .ZN(SubCellInst_LFInst_8_n21) );
  OAI22_X1 SubCellInst_LFInst_9_U11 ( .A1(Output[31]), .A2(Output[28]), .B1(
        SubCellInst_LFInst_9_n27), .B2(Output[29]), .ZN(Feedback[39]) );
  NOR2_X1 SubCellInst_LFInst_9_U10 ( .A1(SubCellInst_LFInst_9_n26), .A2(
        SubCellInst_LFInst_9_n25), .ZN(SubCellInst_LFInst_9_n27) );
  OAI22_X1 SubCellInst_LFInst_9_U9 ( .A1(Output[31]), .A2(Output[28]), .B1(
        SubCellInst_LFInst_9_n24), .B2(SubCellInst_LFInst_9_n23), .ZN(
        Feedback[38]) );
  AOI21_X1 SubCellInst_LFInst_9_U8 ( .B1(Output[28]), .B2(Output[31]), .A(
        Output[30]), .ZN(SubCellInst_LFInst_9_n23) );
  OAI21_X1 SubCellInst_LFInst_9_U7 ( .B1(Output[31]), .B2(
        SubCellInst_LFInst_9_n26), .A(SubCellInst_LFInst_9_n22), .ZN(
        Feedback[37]) );
  OAI21_X1 SubCellInst_LFInst_9_U6 ( .B1(Output[30]), .B2(
        SubCellInst_LFInst_9_n25), .A(Output[28]), .ZN(
        SubCellInst_LFInst_9_n22) );
  INV_X1 SubCellInst_LFInst_9_U5 ( .A(Output[31]), .ZN(
        SubCellInst_LFInst_9_n25) );
  INV_X1 SubCellInst_LFInst_9_U4 ( .A(Output[30]), .ZN(
        SubCellInst_LFInst_9_n26) );
  AOI22_X1 SubCellInst_LFInst_9_U3 ( .A1(Output[31]), .A2(Output[30]), .B1(
        SubCellInst_LFInst_9_n21), .B2(SubCellInst_LFInst_9_n24), .ZN(
        Feedback[36]) );
  INV_X1 SubCellInst_LFInst_9_U2 ( .A(Output[29]), .ZN(
        SubCellInst_LFInst_9_n24) );
  OAI21_X1 SubCellInst_LFInst_9_U1 ( .B1(Output[30]), .B2(Output[31]), .A(
        Output[28]), .ZN(SubCellInst_LFInst_9_n21) );
  OAI22_X1 SubCellInst_LFInst_10_U11 ( .A1(Output[27]), .A2(Output[24]), .B1(
        SubCellInst_LFInst_10_n27), .B2(Output[25]), .ZN(Feedback[43]) );
  NOR2_X1 SubCellInst_LFInst_10_U10 ( .A1(SubCellInst_LFInst_10_n26), .A2(
        SubCellInst_LFInst_10_n25), .ZN(SubCellInst_LFInst_10_n27) );
  OAI22_X1 SubCellInst_LFInst_10_U9 ( .A1(Output[27]), .A2(Output[24]), .B1(
        SubCellInst_LFInst_10_n24), .B2(SubCellInst_LFInst_10_n23), .ZN(
        Feedback[42]) );
  AOI21_X1 SubCellInst_LFInst_10_U8 ( .B1(Output[24]), .B2(Output[27]), .A(
        Output[26]), .ZN(SubCellInst_LFInst_10_n23) );
  OAI21_X1 SubCellInst_LFInst_10_U7 ( .B1(Output[27]), .B2(
        SubCellInst_LFInst_10_n26), .A(SubCellInst_LFInst_10_n22), .ZN(
        Feedback[41]) );
  OAI21_X1 SubCellInst_LFInst_10_U6 ( .B1(Output[26]), .B2(
        SubCellInst_LFInst_10_n25), .A(Output[24]), .ZN(
        SubCellInst_LFInst_10_n22) );
  INV_X1 SubCellInst_LFInst_10_U5 ( .A(Output[27]), .ZN(
        SubCellInst_LFInst_10_n25) );
  INV_X1 SubCellInst_LFInst_10_U4 ( .A(Output[26]), .ZN(
        SubCellInst_LFInst_10_n26) );
  AOI22_X1 SubCellInst_LFInst_10_U3 ( .A1(Output[27]), .A2(Output[26]), .B1(
        SubCellInst_LFInst_10_n21), .B2(SubCellInst_LFInst_10_n24), .ZN(
        Feedback[40]) );
  INV_X1 SubCellInst_LFInst_10_U2 ( .A(Output[25]), .ZN(
        SubCellInst_LFInst_10_n24) );
  OAI21_X1 SubCellInst_LFInst_10_U1 ( .B1(Output[26]), .B2(Output[27]), .A(
        Output[24]), .ZN(SubCellInst_LFInst_10_n21) );
  OAI22_X1 SubCellInst_LFInst_11_U11 ( .A1(Output[23]), .A2(Output[20]), .B1(
        SubCellInst_LFInst_11_n27), .B2(Output[21]), .ZN(Feedback[47]) );
  NOR2_X1 SubCellInst_LFInst_11_U10 ( .A1(SubCellInst_LFInst_11_n26), .A2(
        SubCellInst_LFInst_11_n25), .ZN(SubCellInst_LFInst_11_n27) );
  OAI22_X1 SubCellInst_LFInst_11_U9 ( .A1(Output[23]), .A2(Output[20]), .B1(
        SubCellInst_LFInst_11_n24), .B2(SubCellInst_LFInst_11_n23), .ZN(
        Feedback[46]) );
  AOI21_X1 SubCellInst_LFInst_11_U8 ( .B1(Output[20]), .B2(Output[23]), .A(
        Output[22]), .ZN(SubCellInst_LFInst_11_n23) );
  OAI21_X1 SubCellInst_LFInst_11_U7 ( .B1(Output[23]), .B2(
        SubCellInst_LFInst_11_n26), .A(SubCellInst_LFInst_11_n22), .ZN(
        Feedback[45]) );
  OAI21_X1 SubCellInst_LFInst_11_U6 ( .B1(Output[22]), .B2(
        SubCellInst_LFInst_11_n25), .A(Output[20]), .ZN(
        SubCellInst_LFInst_11_n22) );
  INV_X1 SubCellInst_LFInst_11_U5 ( .A(Output[23]), .ZN(
        SubCellInst_LFInst_11_n25) );
  INV_X1 SubCellInst_LFInst_11_U4 ( .A(Output[22]), .ZN(
        SubCellInst_LFInst_11_n26) );
  AOI22_X1 SubCellInst_LFInst_11_U3 ( .A1(Output[23]), .A2(Output[22]), .B1(
        SubCellInst_LFInst_11_n21), .B2(SubCellInst_LFInst_11_n24), .ZN(
        Feedback[44]) );
  INV_X1 SubCellInst_LFInst_11_U2 ( .A(Output[21]), .ZN(
        SubCellInst_LFInst_11_n24) );
  OAI21_X1 SubCellInst_LFInst_11_U1 ( .B1(Output[22]), .B2(Output[23]), .A(
        Output[20]), .ZN(SubCellInst_LFInst_11_n21) );
  OAI22_X1 SubCellInst_LFInst_12_U11 ( .A1(Output[7]), .A2(Output[4]), .B1(
        SubCellInst_LFInst_12_n27), .B2(Output[5]), .ZN(Feedback[51]) );
  NOR2_X1 SubCellInst_LFInst_12_U10 ( .A1(SubCellInst_LFInst_12_n26), .A2(
        SubCellInst_LFInst_12_n25), .ZN(SubCellInst_LFInst_12_n27) );
  OAI22_X1 SubCellInst_LFInst_12_U9 ( .A1(Output[7]), .A2(Output[4]), .B1(
        SubCellInst_LFInst_12_n24), .B2(SubCellInst_LFInst_12_n23), .ZN(
        Feedback[50]) );
  AOI21_X1 SubCellInst_LFInst_12_U8 ( .B1(Output[4]), .B2(Output[7]), .A(
        Output[6]), .ZN(SubCellInst_LFInst_12_n23) );
  OAI21_X1 SubCellInst_LFInst_12_U7 ( .B1(Output[7]), .B2(
        SubCellInst_LFInst_12_n26), .A(SubCellInst_LFInst_12_n22), .ZN(
        Feedback[49]) );
  OAI21_X1 SubCellInst_LFInst_12_U6 ( .B1(Output[6]), .B2(
        SubCellInst_LFInst_12_n25), .A(Output[4]), .ZN(
        SubCellInst_LFInst_12_n22) );
  INV_X1 SubCellInst_LFInst_12_U5 ( .A(Output[7]), .ZN(
        SubCellInst_LFInst_12_n25) );
  INV_X1 SubCellInst_LFInst_12_U4 ( .A(Output[6]), .ZN(
        SubCellInst_LFInst_12_n26) );
  AOI22_X1 SubCellInst_LFInst_12_U3 ( .A1(Output[7]), .A2(Output[6]), .B1(
        SubCellInst_LFInst_12_n21), .B2(SubCellInst_LFInst_12_n24), .ZN(
        Feedback[48]) );
  INV_X1 SubCellInst_LFInst_12_U2 ( .A(Output[5]), .ZN(
        SubCellInst_LFInst_12_n24) );
  OAI21_X1 SubCellInst_LFInst_12_U1 ( .B1(Output[6]), .B2(Output[7]), .A(
        Output[4]), .ZN(SubCellInst_LFInst_12_n21) );
  OAI22_X1 SubCellInst_LFInst_13_U11 ( .A1(Output[11]), .A2(Output[8]), .B1(
        SubCellInst_LFInst_13_n27), .B2(Output[9]), .ZN(Feedback[55]) );
  NOR2_X1 SubCellInst_LFInst_13_U10 ( .A1(SubCellInst_LFInst_13_n26), .A2(
        SubCellInst_LFInst_13_n25), .ZN(SubCellInst_LFInst_13_n27) );
  OAI22_X1 SubCellInst_LFInst_13_U9 ( .A1(Output[11]), .A2(Output[8]), .B1(
        SubCellInst_LFInst_13_n24), .B2(SubCellInst_LFInst_13_n23), .ZN(
        Feedback[54]) );
  AOI21_X1 SubCellInst_LFInst_13_U8 ( .B1(Output[8]), .B2(Output[11]), .A(
        Output[10]), .ZN(SubCellInst_LFInst_13_n23) );
  OAI21_X1 SubCellInst_LFInst_13_U7 ( .B1(Output[11]), .B2(
        SubCellInst_LFInst_13_n26), .A(SubCellInst_LFInst_13_n22), .ZN(
        Feedback[53]) );
  OAI21_X1 SubCellInst_LFInst_13_U6 ( .B1(Output[10]), .B2(
        SubCellInst_LFInst_13_n25), .A(Output[8]), .ZN(
        SubCellInst_LFInst_13_n22) );
  INV_X1 SubCellInst_LFInst_13_U5 ( .A(Output[11]), .ZN(
        SubCellInst_LFInst_13_n25) );
  INV_X1 SubCellInst_LFInst_13_U4 ( .A(Output[10]), .ZN(
        SubCellInst_LFInst_13_n26) );
  AOI22_X1 SubCellInst_LFInst_13_U3 ( .A1(Output[11]), .A2(Output[10]), .B1(
        SubCellInst_LFInst_13_n21), .B2(SubCellInst_LFInst_13_n24), .ZN(
        Feedback[52]) );
  INV_X1 SubCellInst_LFInst_13_U2 ( .A(Output[9]), .ZN(
        SubCellInst_LFInst_13_n24) );
  OAI21_X1 SubCellInst_LFInst_13_U1 ( .B1(Output[10]), .B2(Output[11]), .A(
        Output[8]), .ZN(SubCellInst_LFInst_13_n21) );
  OAI22_X1 SubCellInst_LFInst_14_U11 ( .A1(Output[15]), .A2(Output[12]), .B1(
        SubCellInst_LFInst_14_n27), .B2(Output[13]), .ZN(Feedback[59]) );
  NOR2_X1 SubCellInst_LFInst_14_U10 ( .A1(SubCellInst_LFInst_14_n26), .A2(
        SubCellInst_LFInst_14_n25), .ZN(SubCellInst_LFInst_14_n27) );
  OAI22_X1 SubCellInst_LFInst_14_U9 ( .A1(Output[15]), .A2(Output[12]), .B1(
        SubCellInst_LFInst_14_n24), .B2(SubCellInst_LFInst_14_n23), .ZN(
        Feedback[58]) );
  AOI21_X1 SubCellInst_LFInst_14_U8 ( .B1(Output[12]), .B2(Output[15]), .A(
        Output[14]), .ZN(SubCellInst_LFInst_14_n23) );
  OAI21_X1 SubCellInst_LFInst_14_U7 ( .B1(Output[15]), .B2(
        SubCellInst_LFInst_14_n26), .A(SubCellInst_LFInst_14_n22), .ZN(
        Feedback[57]) );
  OAI21_X1 SubCellInst_LFInst_14_U6 ( .B1(Output[14]), .B2(
        SubCellInst_LFInst_14_n25), .A(Output[12]), .ZN(
        SubCellInst_LFInst_14_n22) );
  INV_X1 SubCellInst_LFInst_14_U5 ( .A(Output[15]), .ZN(
        SubCellInst_LFInst_14_n25) );
  INV_X1 SubCellInst_LFInst_14_U4 ( .A(Output[14]), .ZN(
        SubCellInst_LFInst_14_n26) );
  AOI22_X1 SubCellInst_LFInst_14_U3 ( .A1(Output[15]), .A2(Output[14]), .B1(
        SubCellInst_LFInst_14_n21), .B2(SubCellInst_LFInst_14_n24), .ZN(
        Feedback[56]) );
  INV_X1 SubCellInst_LFInst_14_U2 ( .A(Output[13]), .ZN(
        SubCellInst_LFInst_14_n24) );
  OAI21_X1 SubCellInst_LFInst_14_U1 ( .B1(Output[14]), .B2(Output[15]), .A(
        Output[12]), .ZN(SubCellInst_LFInst_14_n21) );
  OAI22_X1 SubCellInst_LFInst_15_U11 ( .A1(Output[3]), .A2(Output[0]), .B1(
        SubCellInst_LFInst_15_n27), .B2(Output[1]), .ZN(Feedback[63]) );
  NOR2_X1 SubCellInst_LFInst_15_U10 ( .A1(SubCellInst_LFInst_15_n26), .A2(
        SubCellInst_LFInst_15_n25), .ZN(SubCellInst_LFInst_15_n27) );
  OAI22_X1 SubCellInst_LFInst_15_U9 ( .A1(Output[3]), .A2(Output[0]), .B1(
        SubCellInst_LFInst_15_n24), .B2(SubCellInst_LFInst_15_n23), .ZN(
        Feedback[62]) );
  AOI21_X1 SubCellInst_LFInst_15_U8 ( .B1(Output[0]), .B2(Output[3]), .A(
        Output[2]), .ZN(SubCellInst_LFInst_15_n23) );
  OAI21_X1 SubCellInst_LFInst_15_U7 ( .B1(Output[3]), .B2(
        SubCellInst_LFInst_15_n26), .A(SubCellInst_LFInst_15_n22), .ZN(
        Feedback[61]) );
  OAI21_X1 SubCellInst_LFInst_15_U6 ( .B1(Output[2]), .B2(
        SubCellInst_LFInst_15_n25), .A(Output[0]), .ZN(
        SubCellInst_LFInst_15_n22) );
  INV_X1 SubCellInst_LFInst_15_U5 ( .A(Output[3]), .ZN(
        SubCellInst_LFInst_15_n25) );
  INV_X1 SubCellInst_LFInst_15_U4 ( .A(Output[2]), .ZN(
        SubCellInst_LFInst_15_n26) );
  AOI22_X1 SubCellInst_LFInst_15_U3 ( .A1(Output[3]), .A2(Output[2]), .B1(
        SubCellInst_LFInst_15_n21), .B2(SubCellInst_LFInst_15_n24), .ZN(
        Feedback[60]) );
  INV_X1 SubCellInst_LFInst_15_U2 ( .A(Output[1]), .ZN(
        SubCellInst_LFInst_15_n24) );
  OAI21_X1 SubCellInst_LFInst_15_U1 ( .B1(Output[2]), .B2(Output[3]), .A(
        Output[0]), .ZN(SubCellInst_LFInst_15_n21) );
  BUF_X1 KeyMUX_U3 ( .A(selects_0_), .Z(KeyMUX_n7) );
  BUF_X1 KeyMUX_U2 ( .A(selects_0_), .Z(KeyMUX_n5) );
  BUF_X1 KeyMUX_U1 ( .A(selects_0_), .Z(KeyMUX_n6) );
  MUX2_X1 KeyMUX_MUXInst_0_U1 ( .A(Key[64]), .B(Key[0]), .S(KeyMUX_n5), .Z(
        SelectedKey[0]) );
  MUX2_X1 KeyMUX_MUXInst_1_U1 ( .A(Key[65]), .B(Key[1]), .S(KeyMUX_n5), .Z(
        SelectedKey[1]) );
  MUX2_X1 KeyMUX_MUXInst_2_U1 ( .A(Key[66]), .B(Key[2]), .S(KeyMUX_n5), .Z(
        SelectedKey[2]) );
  MUX2_X1 KeyMUX_MUXInst_3_U1 ( .A(Key[67]), .B(Key[3]), .S(KeyMUX_n5), .Z(
        SelectedKey[3]) );
  MUX2_X1 KeyMUX_MUXInst_4_U1 ( .A(Key[68]), .B(Key[4]), .S(KeyMUX_n5), .Z(
        SelectedKey[4]) );
  MUX2_X1 KeyMUX_MUXInst_5_U1 ( .A(Key[69]), .B(Key[5]), .S(KeyMUX_n5), .Z(
        SelectedKey[5]) );
  MUX2_X1 KeyMUX_MUXInst_6_U1 ( .A(Key[70]), .B(Key[6]), .S(KeyMUX_n5), .Z(
        SelectedKey[6]) );
  MUX2_X1 KeyMUX_MUXInst_7_U1 ( .A(Key[71]), .B(Key[7]), .S(KeyMUX_n5), .Z(
        SelectedKey[7]) );
  MUX2_X1 KeyMUX_MUXInst_8_U1 ( .A(Key[72]), .B(Key[8]), .S(KeyMUX_n5), .Z(
        SelectedKey[8]) );
  MUX2_X1 KeyMUX_MUXInst_9_U1 ( .A(Key[73]), .B(Key[9]), .S(KeyMUX_n5), .Z(
        SelectedKey[9]) );
  MUX2_X1 KeyMUX_MUXInst_10_U1 ( .A(Key[74]), .B(Key[10]), .S(KeyMUX_n5), .Z(
        SelectedKey[10]) );
  MUX2_X1 KeyMUX_MUXInst_11_U1 ( .A(Key[75]), .B(Key[11]), .S(KeyMUX_n5), .Z(
        SelectedKey[11]) );
  MUX2_X1 KeyMUX_MUXInst_12_U1 ( .A(Key[76]), .B(Key[12]), .S(KeyMUX_n6), .Z(
        SelectedKey[12]) );
  MUX2_X1 KeyMUX_MUXInst_13_U1 ( .A(Key[77]), .B(Key[13]), .S(KeyMUX_n6), .Z(
        SelectedKey[13]) );
  MUX2_X1 KeyMUX_MUXInst_14_U1 ( .A(Key[78]), .B(Key[14]), .S(KeyMUX_n6), .Z(
        SelectedKey[14]) );
  MUX2_X1 KeyMUX_MUXInst_15_U1 ( .A(Key[79]), .B(Key[15]), .S(KeyMUX_n6), .Z(
        SelectedKey[15]) );
  MUX2_X1 KeyMUX_MUXInst_16_U1 ( .A(Key[80]), .B(Key[16]), .S(KeyMUX_n6), .Z(
        SelectedKey[16]) );
  MUX2_X1 KeyMUX_MUXInst_17_U1 ( .A(Key[81]), .B(Key[17]), .S(KeyMUX_n6), .Z(
        SelectedKey[17]) );
  MUX2_X1 KeyMUX_MUXInst_18_U1 ( .A(Key[82]), .B(Key[18]), .S(KeyMUX_n6), .Z(
        SelectedKey[18]) );
  MUX2_X1 KeyMUX_MUXInst_19_U1 ( .A(Key[83]), .B(Key[19]), .S(KeyMUX_n6), .Z(
        SelectedKey[19]) );
  MUX2_X1 KeyMUX_MUXInst_20_U1 ( .A(Key[84]), .B(Key[20]), .S(KeyMUX_n6), .Z(
        SelectedKey[20]) );
  MUX2_X1 KeyMUX_MUXInst_21_U1 ( .A(Key[85]), .B(Key[21]), .S(KeyMUX_n6), .Z(
        SelectedKey[21]) );
  MUX2_X1 KeyMUX_MUXInst_22_U1 ( .A(Key[86]), .B(Key[22]), .S(KeyMUX_n6), .Z(
        SelectedKey[22]) );
  MUX2_X1 KeyMUX_MUXInst_23_U1 ( .A(Key[87]), .B(Key[23]), .S(KeyMUX_n6), .Z(
        SelectedKey[23]) );
  MUX2_X1 KeyMUX_MUXInst_24_U1 ( .A(Key[88]), .B(Key[24]), .S(KeyMUX_n7), .Z(
        SelectedKey[24]) );
  MUX2_X1 KeyMUX_MUXInst_25_U1 ( .A(Key[89]), .B(Key[25]), .S(KeyMUX_n7), .Z(
        SelectedKey[25]) );
  MUX2_X1 KeyMUX_MUXInst_26_U1 ( .A(Key[90]), .B(Key[26]), .S(KeyMUX_n7), .Z(
        SelectedKey[26]) );
  MUX2_X1 KeyMUX_MUXInst_27_U1 ( .A(Key[91]), .B(Key[27]), .S(KeyMUX_n7), .Z(
        SelectedKey[27]) );
  MUX2_X1 KeyMUX_MUXInst_28_U1 ( .A(Key[92]), .B(Key[28]), .S(KeyMUX_n7), .Z(
        SelectedKey[28]) );
  MUX2_X1 KeyMUX_MUXInst_29_U1 ( .A(Key[93]), .B(Key[29]), .S(KeyMUX_n7), .Z(
        SelectedKey[29]) );
  MUX2_X1 KeyMUX_MUXInst_30_U1 ( .A(Key[94]), .B(Key[30]), .S(KeyMUX_n7), .Z(
        SelectedKey[30]) );
  MUX2_X1 KeyMUX_MUXInst_31_U1 ( .A(Key[95]), .B(Key[31]), .S(KeyMUX_n7), .Z(
        SelectedKey[31]) );
  MUX2_X1 KeyMUX_MUXInst_32_U1 ( .A(Key[96]), .B(Key[32]), .S(KeyMUX_n7), .Z(
        SelectedKey[32]) );
  MUX2_X1 KeyMUX_MUXInst_33_U1 ( .A(Key[97]), .B(Key[33]), .S(KeyMUX_n7), .Z(
        SelectedKey[33]) );
  MUX2_X1 KeyMUX_MUXInst_34_U1 ( .A(Key[98]), .B(Key[34]), .S(KeyMUX_n7), .Z(
        SelectedKey[34]) );
  MUX2_X1 KeyMUX_MUXInst_35_U1 ( .A(Key[99]), .B(Key[35]), .S(KeyMUX_n7), .Z(
        SelectedKey[35]) );
  MUX2_X1 KeyMUX_MUXInst_36_U1 ( .A(Key[100]), .B(Key[36]), .S(KeyMUX_n7), .Z(
        SelectedKey[36]) );
  MUX2_X1 KeyMUX_MUXInst_37_U1 ( .A(Key[101]), .B(Key[37]), .S(KeyMUX_n7), .Z(
        SelectedKey[37]) );
  MUX2_X1 KeyMUX_MUXInst_38_U1 ( .A(Key[102]), .B(Key[38]), .S(KeyMUX_n7), .Z(
        SelectedKey[38]) );
  MUX2_X1 KeyMUX_MUXInst_39_U1 ( .A(Key[103]), .B(Key[39]), .S(KeyMUX_n7), .Z(
        SelectedKey[39]) );
  MUX2_X1 KeyMUX_MUXInst_40_U1 ( .A(Key[104]), .B(Key[40]), .S(selects_0_), 
        .Z(SelectedKey[40]) );
  MUX2_X1 KeyMUX_MUXInst_41_U1 ( .A(Key[105]), .B(Key[41]), .S(KeyMUX_n7), .Z(
        SelectedKey[41]) );
  MUX2_X1 KeyMUX_MUXInst_42_U1 ( .A(Key[106]), .B(Key[42]), .S(selects_0_), 
        .Z(SelectedKey[42]) );
  MUX2_X1 KeyMUX_MUXInst_43_U1 ( .A(Key[107]), .B(Key[43]), .S(KeyMUX_n7), .Z(
        SelectedKey[43]) );
  MUX2_X1 KeyMUX_MUXInst_44_U1 ( .A(Key[108]), .B(Key[44]), .S(selects_0_), 
        .Z(SelectedKey[44]) );
  MUX2_X1 KeyMUX_MUXInst_45_U1 ( .A(Key[109]), .B(Key[45]), .S(KeyMUX_n7), .Z(
        SelectedKey[45]) );
  MUX2_X1 KeyMUX_MUXInst_46_U1 ( .A(Key[110]), .B(Key[46]), .S(selects_0_), 
        .Z(SelectedKey[46]) );
  MUX2_X1 KeyMUX_MUXInst_47_U1 ( .A(Key[111]), .B(Key[47]), .S(selects_0_), 
        .Z(SelectedKey[47]) );
  MUX2_X1 KeyMUX_MUXInst_48_U1 ( .A(Key[112]), .B(Key[48]), .S(KeyMUX_n6), .Z(
        SelectedKey[48]) );
  MUX2_X1 KeyMUX_MUXInst_49_U1 ( .A(Key[113]), .B(Key[49]), .S(KeyMUX_n5), .Z(
        SelectedKey[49]) );
  MUX2_X1 KeyMUX_MUXInst_50_U1 ( .A(Key[114]), .B(Key[50]), .S(KeyMUX_n6), .Z(
        SelectedKey[50]) );
  MUX2_X1 KeyMUX_MUXInst_51_U1 ( .A(Key[115]), .B(Key[51]), .S(KeyMUX_n5), .Z(
        SelectedKey[51]) );
  MUX2_X1 KeyMUX_MUXInst_52_U1 ( .A(Key[116]), .B(Key[52]), .S(KeyMUX_n6), .Z(
        SelectedKey[52]) );
  MUX2_X1 KeyMUX_MUXInst_53_U1 ( .A(Key[117]), .B(Key[53]), .S(KeyMUX_n5), .Z(
        SelectedKey[53]) );
  MUX2_X1 KeyMUX_MUXInst_54_U1 ( .A(Key[118]), .B(Key[54]), .S(KeyMUX_n6), .Z(
        SelectedKey[54]) );
  MUX2_X1 KeyMUX_MUXInst_55_U1 ( .A(Key[119]), .B(Key[55]), .S(KeyMUX_n5), .Z(
        SelectedKey[55]) );
  MUX2_X1 KeyMUX_MUXInst_56_U1 ( .A(Key[120]), .B(Key[56]), .S(KeyMUX_n6), .Z(
        SelectedKey[56]) );
  MUX2_X1 KeyMUX_MUXInst_57_U1 ( .A(Key[121]), .B(Key[57]), .S(KeyMUX_n5), .Z(
        SelectedKey[57]) );
  MUX2_X1 KeyMUX_MUXInst_58_U1 ( .A(Key[122]), .B(Key[58]), .S(KeyMUX_n6), .Z(
        SelectedKey[58]) );
  MUX2_X1 KeyMUX_MUXInst_59_U1 ( .A(Key[123]), .B(Key[59]), .S(KeyMUX_n5), .Z(
        SelectedKey[59]) );
  MUX2_X1 KeyMUX_MUXInst_60_U1 ( .A(Key[124]), .B(Key[60]), .S(KeyMUX_n6), .Z(
        SelectedKey[60]) );
  MUX2_X1 KeyMUX_MUXInst_61_U1 ( .A(Key[125]), .B(Key[61]), .S(KeyMUX_n7), .Z(
        SelectedKey[61]) );
  MUX2_X1 KeyMUX_MUXInst_62_U1 ( .A(Key[126]), .B(Key[62]), .S(KeyMUX_n6), .Z(
        SelectedKey[62]) );
  MUX2_X1 KeyMUX_MUXInst_63_U1 ( .A(Key[127]), .B(Key[63]), .S(KeyMUX_n5), .Z(
        SelectedKey[63]) );
  OR2_X1 FSMMUX_MUXInst_0_U1 ( .A1(FSMReg[0]), .A2(rst), .ZN(RoundConstant_0)
         );
  NOR2_X1 FSMMUX_MUXInst_1_U2 ( .A1(rst), .A2(FSMMUX_MUXInst_1_n4), .ZN(
        FSMUpdate[0]) );
  INV_X1 FSMMUX_MUXInst_1_U1 ( .A(FSMReg[1]), .ZN(FSMMUX_MUXInst_1_n4) );
  NOR2_X1 FSMMUX_MUXInst_2_U2 ( .A1(rst), .A2(FSMMUX_MUXInst_2_n4), .ZN(
        FSMUpdate[1]) );
  INV_X1 FSMMUX_MUXInst_2_U1 ( .A(FSMReg[2]), .ZN(FSMMUX_MUXInst_2_n4) );
  OR2_X1 FSMMUX_MUXInst_3_U1 ( .A1(FSMReg[3]), .A2(rst), .ZN(RoundConstant_4_)
         );
  NOR2_X1 FSMMUX_MUXInst_4_U2 ( .A1(rst), .A2(FSMMUX_MUXInst_4_n4), .ZN(
        FSMUpdate[3]) );
  INV_X1 FSMMUX_MUXInst_4_U1 ( .A(FSMReg[4]), .ZN(FSMMUX_MUXInst_4_n4) );
  NOR2_X1 FSMMUX_MUXInst_5_U2 ( .A1(rst), .A2(FSMMUX_MUXInst_5_n4), .ZN(
        FSMUpdate[4]) );
  INV_X1 FSMMUX_MUXInst_5_U1 ( .A(FSMReg[5]), .ZN(FSMMUX_MUXInst_5_n4) );
  NOR2_X1 FSMMUX_MUXInst_6_U2 ( .A1(rst), .A2(FSMMUX_MUXInst_6_n4), .ZN(
        FSMUpdate[5]) );
  INV_X1 FSMMUX_MUXInst_6_U1 ( .A(FSMReg[6]), .ZN(FSMMUX_MUXInst_6_n4) );
  XOR2_X1 FSMUpdateInst_U2 ( .A(RoundConstant_4_), .B(FSMUpdate[3]), .Z(
        FSMUpdate[6]) );
  XOR2_X1 FSMUpdateInst_U1 ( .A(FSMUpdate[0]), .B(RoundConstant_0), .Z(
        FSMUpdate[2]) );
  DFF_X1 FSMRegInst_s_current_state_reg_0_ ( .D(FSMUpdate[0]), .CK(clk), .Q(
        FSMReg[0]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_1_ ( .D(FSMUpdate[1]), .CK(clk), .Q(
        FSMReg[1]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_2_ ( .D(FSMUpdate[2]), .CK(clk), .Q(
        FSMReg[2]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_3_ ( .D(FSMUpdate[3]), .CK(clk), .Q(
        FSMReg[3]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_4_ ( .D(FSMUpdate[4]), .CK(clk), .Q(
        FSMReg[4]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_5_ ( .D(FSMUpdate[5]), .CK(clk), .Q(
        FSMReg[5]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_6_ ( .D(FSMUpdate[6]), .CK(clk), .Q(
        FSMReg[6]), .QN() );
  AND4_X1 FSMSignalsInst_U2 ( .A1(RoundConstant_0), .A2(FSMUpdate[1]), .A3(
        FSMUpdate[5]), .A4(FSMSignalsInst_n1), .ZN(done) );
  NOR4_X1 FSMSignalsInst_U1 ( .A1(FSMUpdate[0]), .A2(RoundConstant_4_), .A3(
        FSMUpdate[3]), .A4(FSMUpdate[4]), .ZN(FSMSignalsInst_n1) );
  MUX2_X1 selectsMUX_MUXInst_0_U1 ( .A(selectsReg_0_), .B(1'b0), .S(rst), 
        .Z(selects_0_) );
  INV_X1 selectsUpdateInst_U1 ( .A(selects_0_), .ZN(selectsNext_0_) );
  DFF_X1 selectsRegInst_s_current_state_reg_0_ ( .D(selectsNext_0_), .CK(clk), 
        .Q(selectsReg_0_), .QN() );
endmodule

