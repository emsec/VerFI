

module Cipher ( clk, rst, EncDec, Input, Key, Tweak, Output, done );
  input [63:0] Input;
  input [127:0] Key;
  input [63:0] Tweak;
  output [63:0] Output;
  input clk, rst, EncDec;
  output done;
  wire   RoundConstant_4_, RoundConstant_0, N3, N4, N5, N6, N7,
         MCInst_XOR_r0_Inst_0_n2, MCInst_XOR_r0_Inst_0_n1,
         MCInst_XOR_r1_Inst_0_n1, MCInst_XOR_r0_Inst_1_n2,
         MCInst_XOR_r0_Inst_1_n1, MCInst_XOR_r1_Inst_1_n1,
         MCInst_XOR_r0_Inst_2_n2, MCInst_XOR_r0_Inst_2_n1,
         MCInst_XOR_r1_Inst_2_n1, MCInst_XOR_r0_Inst_3_n2,
         MCInst_XOR_r0_Inst_3_n1, MCInst_XOR_r1_Inst_3_n1,
         MCInst_XOR_r0_Inst_4_n2, MCInst_XOR_r0_Inst_4_n1,
         MCInst_XOR_r1_Inst_4_n1, MCInst_XOR_r0_Inst_5_n2,
         MCInst_XOR_r0_Inst_5_n1, MCInst_XOR_r1_Inst_5_n1,
         MCInst_XOR_r0_Inst_6_n2, MCInst_XOR_r0_Inst_6_n1,
         MCInst_XOR_r1_Inst_6_n1, MCInst_XOR_r0_Inst_7_n2,
         MCInst_XOR_r0_Inst_7_n1, MCInst_XOR_r1_Inst_7_n1,
         MCInst_XOR_r0_Inst_8_n2, MCInst_XOR_r0_Inst_8_n1,
         MCInst_XOR_r1_Inst_8_n1, MCInst_XOR_r0_Inst_9_n2,
         MCInst_XOR_r0_Inst_9_n1, MCInst_XOR_r1_Inst_9_n1,
         MCInst_XOR_r0_Inst_10_n2, MCInst_XOR_r0_Inst_10_n1,
         MCInst_XOR_r1_Inst_10_n1, MCInst_XOR_r0_Inst_11_n2,
         MCInst_XOR_r0_Inst_11_n1, MCInst_XOR_r1_Inst_11_n1,
         MCInst_XOR_r0_Inst_12_n2, MCInst_XOR_r0_Inst_12_n1,
         MCInst_XOR_r1_Inst_12_n1, MCInst_XOR_r0_Inst_13_n2,
         MCInst_XOR_r0_Inst_13_n1, MCInst_XOR_r1_Inst_13_n1,
         MCInst_XOR_r0_Inst_14_n2, MCInst_XOR_r0_Inst_14_n1,
         MCInst_XOR_r1_Inst_14_n1, MCInst_XOR_r0_Inst_15_n2,
         MCInst_XOR_r0_Inst_15_n1, MCInst_XOR_r1_Inst_15_n1,
         AddKeyXOR1_XORInst_0_0_n1, AddKeyXOR1_XORInst_0_1_n1,
         AddKeyXOR1_XORInst_0_2_n1, AddKeyXOR1_XORInst_0_3_n1,
         AddKeyXOR1_XORInst_1_0_n1, AddKeyXOR1_XORInst_1_1_n1,
         AddKeyXOR1_XORInst_1_2_n1, AddKeyXOR1_XORInst_1_3_n1,
         AddKeyXOR1_XORInst_2_0_n1, AddKeyXOR1_XORInst_2_1_n1,
         AddKeyXOR1_XORInst_2_2_n1, AddKeyXOR1_XORInst_2_3_n1,
         AddKeyXOR1_XORInst_3_0_n1, AddKeyXOR1_XORInst_3_1_n1,
         AddKeyXOR1_XORInst_3_2_n1, AddKeyXOR1_XORInst_3_3_n1,
         AddKeyConstXOR_XORInst_0_0_n2, AddKeyConstXOR_XORInst_0_0_n1,
         AddKeyConstXOR_XORInst_0_1_n2, AddKeyConstXOR_XORInst_0_1_n1,
         AddKeyConstXOR_XORInst_0_2_n2, AddKeyConstXOR_XORInst_0_2_n1,
         AddKeyConstXOR_XORInst_0_3_n2, AddKeyConstXOR_XORInst_0_3_n1,
         AddKeyConstXOR_XORInst_1_0_n2, AddKeyConstXOR_XORInst_1_0_n1,
         AddKeyConstXOR_XORInst_1_1_n2, AddKeyConstXOR_XORInst_1_1_n1,
         AddKeyConstXOR_XORInst_1_2_n2, AddKeyConstXOR_XORInst_1_2_n1,
         AddKeyConstXOR_XORInst_1_3_n2, AddKeyConstXOR_XORInst_1_3_n1,
         AddKeyXOR2_XORInst_0_0_n1, AddKeyXOR2_XORInst_0_1_n1,
         AddKeyXOR2_XORInst_0_2_n1, AddKeyXOR2_XORInst_0_3_n1,
         AddKeyXOR2_XORInst_1_0_n1, AddKeyXOR2_XORInst_1_1_n1,
         AddKeyXOR2_XORInst_1_2_n1, AddKeyXOR2_XORInst_1_3_n1,
         AddKeyXOR2_XORInst_2_0_n1, AddKeyXOR2_XORInst_2_1_n1,
         AddKeyXOR2_XORInst_2_2_n1, AddKeyXOR2_XORInst_2_3_n1,
         AddKeyXOR2_XORInst_3_0_n1, AddKeyXOR2_XORInst_3_1_n1,
         AddKeyXOR2_XORInst_3_2_n1, AddKeyXOR2_XORInst_3_3_n1,
         AddKeyXOR2_XORInst_4_0_n1, AddKeyXOR2_XORInst_4_1_n1,
         AddKeyXOR2_XORInst_4_2_n1, AddKeyXOR2_XORInst_4_3_n1,
         AddKeyXOR2_XORInst_5_0_n1, AddKeyXOR2_XORInst_5_1_n1,
         AddKeyXOR2_XORInst_5_2_n1, AddKeyXOR2_XORInst_5_3_n1,
         AddKeyXOR2_XORInst_6_0_n1, AddKeyXOR2_XORInst_6_1_n1,
         AddKeyXOR2_XORInst_6_2_n1, AddKeyXOR2_XORInst_6_3_n1,
         AddKeyXOR2_XORInst_7_0_n1, AddKeyXOR2_XORInst_7_1_n1,
         AddKeyXOR2_XORInst_7_2_n1, AddKeyXOR2_XORInst_7_3_n1,
         AddKeyXOR2_XORInst_8_0_n1, AddKeyXOR2_XORInst_8_1_n1,
         AddKeyXOR2_XORInst_8_2_n1, AddKeyXOR2_XORInst_8_3_n1,
         AddKeyXOR2_XORInst_9_0_n1, AddKeyXOR2_XORInst_9_1_n1,
         AddKeyXOR2_XORInst_9_2_n1, AddKeyXOR2_XORInst_9_3_n1,
         SubCellInst_LFInst_0_LFInst_0_n1, SubCellInst_LFInst_0_LFInst_1_n2,
         SubCellInst_LFInst_0_LFInst_1_n1, SubCellInst_LFInst_0_LFInst_2_n1,
         SubCellInst_LFInst_1_LFInst_0_n1, SubCellInst_LFInst_1_LFInst_1_n2,
         SubCellInst_LFInst_1_LFInst_1_n1, SubCellInst_LFInst_1_LFInst_2_n1,
         SubCellInst_LFInst_2_LFInst_0_n1, SubCellInst_LFInst_2_LFInst_1_n2,
         SubCellInst_LFInst_2_LFInst_1_n1, SubCellInst_LFInst_2_LFInst_2_n1,
         SubCellInst_LFInst_3_LFInst_0_n1, SubCellInst_LFInst_3_LFInst_1_n2,
         SubCellInst_LFInst_3_LFInst_1_n1, SubCellInst_LFInst_3_LFInst_2_n1,
         SubCellInst_LFInst_4_LFInst_0_n1, SubCellInst_LFInst_4_LFInst_1_n2,
         SubCellInst_LFInst_4_LFInst_1_n1, SubCellInst_LFInst_4_LFInst_2_n1,
         SubCellInst_LFInst_5_LFInst_0_n1, SubCellInst_LFInst_5_LFInst_1_n2,
         SubCellInst_LFInst_5_LFInst_1_n1, SubCellInst_LFInst_5_LFInst_2_n1,
         SubCellInst_LFInst_6_LFInst_0_n1, SubCellInst_LFInst_6_LFInst_1_n2,
         SubCellInst_LFInst_6_LFInst_1_n1, SubCellInst_LFInst_6_LFInst_2_n1,
         SubCellInst_LFInst_7_LFInst_0_n1, SubCellInst_LFInst_7_LFInst_1_n2,
         SubCellInst_LFInst_7_LFInst_1_n1, SubCellInst_LFInst_7_LFInst_2_n1,
         SubCellInst_LFInst_8_LFInst_0_n1, SubCellInst_LFInst_8_LFInst_1_n2,
         SubCellInst_LFInst_8_LFInst_1_n1, SubCellInst_LFInst_8_LFInst_2_n1,
         SubCellInst_LFInst_9_LFInst_0_n1, SubCellInst_LFInst_9_LFInst_1_n2,
         SubCellInst_LFInst_9_LFInst_1_n1, SubCellInst_LFInst_9_LFInst_2_n1,
         SubCellInst_LFInst_10_LFInst_0_n1, SubCellInst_LFInst_10_LFInst_1_n2,
         SubCellInst_LFInst_10_LFInst_1_n1, SubCellInst_LFInst_10_LFInst_2_n1,
         SubCellInst_LFInst_11_LFInst_0_n1, SubCellInst_LFInst_11_LFInst_1_n2,
         SubCellInst_LFInst_11_LFInst_1_n1, SubCellInst_LFInst_11_LFInst_2_n1,
         SubCellInst_LFInst_12_LFInst_0_n1, SubCellInst_LFInst_12_LFInst_1_n2,
         SubCellInst_LFInst_12_LFInst_1_n1, SubCellInst_LFInst_12_LFInst_2_n1,
         SubCellInst_LFInst_13_LFInst_0_n1, SubCellInst_LFInst_13_LFInst_1_n2,
         SubCellInst_LFInst_13_LFInst_1_n1, SubCellInst_LFInst_13_LFInst_2_n1,
         SubCellInst_LFInst_14_LFInst_0_n1, SubCellInst_LFInst_14_LFInst_1_n2,
         SubCellInst_LFInst_14_LFInst_1_n1, SubCellInst_LFInst_14_LFInst_2_n1,
         SubCellInst_LFInst_15_LFInst_0_n1, SubCellInst_LFInst_15_LFInst_1_n2,
         SubCellInst_LFInst_15_LFInst_1_n1, SubCellInst_LFInst_15_LFInst_2_n1,
         Red_PlaintextInst_LFInst_0_LFInst_0_n1,
         Red_PlaintextInst_LFInst_0_LFInst_1_n1,
         Red_PlaintextInst_LFInst_0_LFInst_2_n1,
         Red_PlaintextInst_LFInst_1_LFInst_0_n1,
         Red_PlaintextInst_LFInst_1_LFInst_1_n1,
         Red_PlaintextInst_LFInst_1_LFInst_2_n1,
         Red_PlaintextInst_LFInst_2_LFInst_0_n1,
         Red_PlaintextInst_LFInst_2_LFInst_1_n1,
         Red_PlaintextInst_LFInst_2_LFInst_2_n1,
         Red_PlaintextInst_LFInst_3_LFInst_0_n1,
         Red_PlaintextInst_LFInst_3_LFInst_1_n1,
         Red_PlaintextInst_LFInst_3_LFInst_2_n1,
         Red_PlaintextInst_LFInst_4_LFInst_0_n1,
         Red_PlaintextInst_LFInst_4_LFInst_1_n1,
         Red_PlaintextInst_LFInst_4_LFInst_2_n1,
         Red_PlaintextInst_LFInst_5_LFInst_0_n1,
         Red_PlaintextInst_LFInst_5_LFInst_1_n1,
         Red_PlaintextInst_LFInst_5_LFInst_2_n1,
         Red_PlaintextInst_LFInst_6_LFInst_0_n1,
         Red_PlaintextInst_LFInst_6_LFInst_1_n1,
         Red_PlaintextInst_LFInst_6_LFInst_2_n1,
         Red_PlaintextInst_LFInst_7_LFInst_0_n1,
         Red_PlaintextInst_LFInst_7_LFInst_1_n1,
         Red_PlaintextInst_LFInst_7_LFInst_2_n1,
         Red_PlaintextInst_LFInst_8_LFInst_0_n1,
         Red_PlaintextInst_LFInst_8_LFInst_1_n1,
         Red_PlaintextInst_LFInst_8_LFInst_2_n1,
         Red_PlaintextInst_LFInst_9_LFInst_0_n1,
         Red_PlaintextInst_LFInst_9_LFInst_1_n1,
         Red_PlaintextInst_LFInst_9_LFInst_2_n1,
         Red_PlaintextInst_LFInst_10_LFInst_0_n1,
         Red_PlaintextInst_LFInst_10_LFInst_1_n1,
         Red_PlaintextInst_LFInst_10_LFInst_2_n1,
         Red_PlaintextInst_LFInst_11_LFInst_0_n1,
         Red_PlaintextInst_LFInst_11_LFInst_1_n1,
         Red_PlaintextInst_LFInst_11_LFInst_2_n1,
         Red_PlaintextInst_LFInst_12_LFInst_0_n1,
         Red_PlaintextInst_LFInst_12_LFInst_1_n1,
         Red_PlaintextInst_LFInst_12_LFInst_2_n1,
         Red_PlaintextInst_LFInst_13_LFInst_0_n1,
         Red_PlaintextInst_LFInst_13_LFInst_1_n1,
         Red_PlaintextInst_LFInst_13_LFInst_2_n1,
         Red_PlaintextInst_LFInst_14_LFInst_0_n1,
         Red_PlaintextInst_LFInst_14_LFInst_1_n1,
         Red_PlaintextInst_LFInst_14_LFInst_2_n1,
         Red_PlaintextInst_LFInst_15_LFInst_0_n1,
         Red_PlaintextInst_LFInst_15_LFInst_1_n1,
         Red_PlaintextInst_LFInst_15_LFInst_2_n1, Red_MCInst_XOR_r0_Inst_0_n2,
         Red_MCInst_XOR_r0_Inst_0_n1, Red_MCInst_XOR_r1_Inst_0_n1,
         Red_MCInst_XOR_r0_Inst_1_n2, Red_MCInst_XOR_r0_Inst_1_n1,
         Red_MCInst_XOR_r1_Inst_1_n1, Red_MCInst_XOR_r0_Inst_2_n2,
         Red_MCInst_XOR_r0_Inst_2_n1, Red_MCInst_XOR_r1_Inst_2_n1,
         Red_MCInst_XOR_r0_Inst_3_n2, Red_MCInst_XOR_r0_Inst_3_n1,
         Red_MCInst_XOR_r1_Inst_3_n1, Red_MCInst_XOR_r0_Inst_4_n2,
         Red_MCInst_XOR_r0_Inst_4_n1, Red_MCInst_XOR_r1_Inst_4_n1,
         Red_MCInst_XOR_r0_Inst_5_n2, Red_MCInst_XOR_r0_Inst_5_n1,
         Red_MCInst_XOR_r1_Inst_5_n1, Red_MCInst_XOR_r0_Inst_6_n2,
         Red_MCInst_XOR_r0_Inst_6_n1, Red_MCInst_XOR_r1_Inst_6_n1,
         Red_MCInst_XOR_r0_Inst_7_n2, Red_MCInst_XOR_r0_Inst_7_n1,
         Red_MCInst_XOR_r1_Inst_7_n1, Red_MCInst_XOR_r0_Inst_8_n2,
         Red_MCInst_XOR_r0_Inst_8_n1, Red_MCInst_XOR_r1_Inst_8_n1,
         Red_MCInst_XOR_r0_Inst_9_n2, Red_MCInst_XOR_r0_Inst_9_n1,
         Red_MCInst_XOR_r1_Inst_9_n1, Red_MCInst_XOR_r0_Inst_10_n2,
         Red_MCInst_XOR_r0_Inst_10_n1, Red_MCInst_XOR_r1_Inst_10_n1,
         Red_MCInst_XOR_r0_Inst_11_n2, Red_MCInst_XOR_r0_Inst_11_n1,
         Red_MCInst_XOR_r1_Inst_11_n1, Red_AddKeyXOR1_XORInst_0_0_n1,
         Red_AddKeyXOR1_XORInst_0_1_n1, Red_AddKeyXOR1_XORInst_0_2_n1,
         Red_AddKeyXOR1_XORInst_1_0_n1, Red_AddKeyXOR1_XORInst_1_1_n1,
         Red_AddKeyXOR1_XORInst_1_2_n1, Red_AddKeyXOR1_XORInst_2_0_n1,
         Red_AddKeyXOR1_XORInst_2_1_n1, Red_AddKeyXOR1_XORInst_2_2_n1,
         Red_AddKeyXOR1_XORInst_3_0_n1, Red_AddKeyXOR1_XORInst_3_1_n1,
         Red_AddKeyXOR1_XORInst_3_2_n1, Red_AddKeyConstXOR_XORInst_0_0_n2,
         Red_AddKeyConstXOR_XORInst_0_0_n1, Red_AddKeyConstXOR_XORInst_0_1_n2,
         Red_AddKeyConstXOR_XORInst_0_1_n1, Red_AddKeyConstXOR_XORInst_0_2_n2,
         Red_AddKeyConstXOR_XORInst_0_2_n1, Red_AddKeyConstXOR_XORInst_1_0_n2,
         Red_AddKeyConstXOR_XORInst_1_0_n1, Red_AddKeyConstXOR_XORInst_1_1_n2,
         Red_AddKeyConstXOR_XORInst_1_1_n1, Red_AddKeyConstXOR_XORInst_1_2_n2,
         Red_AddKeyConstXOR_XORInst_1_2_n1, Red_AddKeyXOR2_XORInst_0_0_n1,
         Red_AddKeyXOR2_XORInst_0_1_n1, Red_AddKeyXOR2_XORInst_0_2_n1,
         Red_AddKeyXOR2_XORInst_1_0_n1, Red_AddKeyXOR2_XORInst_1_1_n1,
         Red_AddKeyXOR2_XORInst_1_2_n1, Red_AddKeyXOR2_XORInst_2_0_n1,
         Red_AddKeyXOR2_XORInst_2_1_n1, Red_AddKeyXOR2_XORInst_2_2_n1,
         Red_AddKeyXOR2_XORInst_3_0_n1, Red_AddKeyXOR2_XORInst_3_1_n1,
         Red_AddKeyXOR2_XORInst_3_2_n1, Red_AddKeyXOR2_XORInst_4_0_n1,
         Red_AddKeyXOR2_XORInst_4_1_n1, Red_AddKeyXOR2_XORInst_4_2_n1,
         Red_AddKeyXOR2_XORInst_5_0_n1, Red_AddKeyXOR2_XORInst_5_1_n1,
         Red_AddKeyXOR2_XORInst_5_2_n1, Red_AddKeyXOR2_XORInst_6_0_n1,
         Red_AddKeyXOR2_XORInst_6_1_n1, Red_AddKeyXOR2_XORInst_6_2_n1,
         Red_AddKeyXOR2_XORInst_7_0_n1, Red_AddKeyXOR2_XORInst_7_1_n1,
         Red_AddKeyXOR2_XORInst_7_2_n1, Red_AddKeyXOR2_XORInst_8_0_n1,
         Red_AddKeyXOR2_XORInst_8_1_n1, Red_AddKeyXOR2_XORInst_8_2_n1,
         Red_AddKeyXOR2_XORInst_9_0_n1, Red_AddKeyXOR2_XORInst_9_1_n1,
         Red_AddKeyXOR2_XORInst_9_2_n1, Red_SubCellInst_LFInst_0_LFInst_0_n2,
         Red_SubCellInst_LFInst_0_LFInst_0_n1,
         Red_SubCellInst_LFInst_0_LFInst_1_n4,
         Red_SubCellInst_LFInst_0_LFInst_1_n3,
         Red_SubCellInst_LFInst_0_LFInst_1_n2,
         Red_SubCellInst_LFInst_0_LFInst_1_n1,
         Red_SubCellInst_LFInst_0_LFInst_2_n6,
         Red_SubCellInst_LFInst_0_LFInst_2_n5,
         Red_SubCellInst_LFInst_0_LFInst_2_n4,
         Red_SubCellInst_LFInst_0_LFInst_2_n3,
         Red_SubCellInst_LFInst_0_LFInst_2_n2,
         Red_SubCellInst_LFInst_0_LFInst_2_n1,
         Red_SubCellInst_LFInst_1_LFInst_0_n2,
         Red_SubCellInst_LFInst_1_LFInst_0_n1,
         Red_SubCellInst_LFInst_1_LFInst_1_n4,
         Red_SubCellInst_LFInst_1_LFInst_1_n3,
         Red_SubCellInst_LFInst_1_LFInst_1_n2,
         Red_SubCellInst_LFInst_1_LFInst_1_n1,
         Red_SubCellInst_LFInst_1_LFInst_2_n6,
         Red_SubCellInst_LFInst_1_LFInst_2_n5,
         Red_SubCellInst_LFInst_1_LFInst_2_n4,
         Red_SubCellInst_LFInst_1_LFInst_2_n3,
         Red_SubCellInst_LFInst_1_LFInst_2_n2,
         Red_SubCellInst_LFInst_1_LFInst_2_n1,
         Red_SubCellInst_LFInst_2_LFInst_0_n2,
         Red_SubCellInst_LFInst_2_LFInst_0_n1,
         Red_SubCellInst_LFInst_2_LFInst_1_n4,
         Red_SubCellInst_LFInst_2_LFInst_1_n3,
         Red_SubCellInst_LFInst_2_LFInst_1_n2,
         Red_SubCellInst_LFInst_2_LFInst_1_n1,
         Red_SubCellInst_LFInst_2_LFInst_2_n6,
         Red_SubCellInst_LFInst_2_LFInst_2_n5,
         Red_SubCellInst_LFInst_2_LFInst_2_n4,
         Red_SubCellInst_LFInst_2_LFInst_2_n3,
         Red_SubCellInst_LFInst_2_LFInst_2_n2,
         Red_SubCellInst_LFInst_2_LFInst_2_n1,
         Red_SubCellInst_LFInst_3_LFInst_0_n2,
         Red_SubCellInst_LFInst_3_LFInst_0_n1,
         Red_SubCellInst_LFInst_3_LFInst_1_n4,
         Red_SubCellInst_LFInst_3_LFInst_1_n3,
         Red_SubCellInst_LFInst_3_LFInst_1_n2,
         Red_SubCellInst_LFInst_3_LFInst_1_n1,
         Red_SubCellInst_LFInst_3_LFInst_2_n6,
         Red_SubCellInst_LFInst_3_LFInst_2_n5,
         Red_SubCellInst_LFInst_3_LFInst_2_n4,
         Red_SubCellInst_LFInst_3_LFInst_2_n3,
         Red_SubCellInst_LFInst_3_LFInst_2_n2,
         Red_SubCellInst_LFInst_3_LFInst_2_n1,
         Red_SubCellInst_LFInst_4_LFInst_0_n2,
         Red_SubCellInst_LFInst_4_LFInst_0_n1,
         Red_SubCellInst_LFInst_4_LFInst_1_n4,
         Red_SubCellInst_LFInst_4_LFInst_1_n3,
         Red_SubCellInst_LFInst_4_LFInst_1_n2,
         Red_SubCellInst_LFInst_4_LFInst_1_n1,
         Red_SubCellInst_LFInst_4_LFInst_2_n6,
         Red_SubCellInst_LFInst_4_LFInst_2_n5,
         Red_SubCellInst_LFInst_4_LFInst_2_n4,
         Red_SubCellInst_LFInst_4_LFInst_2_n3,
         Red_SubCellInst_LFInst_4_LFInst_2_n2,
         Red_SubCellInst_LFInst_4_LFInst_2_n1,
         Red_SubCellInst_LFInst_5_LFInst_0_n2,
         Red_SubCellInst_LFInst_5_LFInst_0_n1,
         Red_SubCellInst_LFInst_5_LFInst_1_n4,
         Red_SubCellInst_LFInst_5_LFInst_1_n3,
         Red_SubCellInst_LFInst_5_LFInst_1_n2,
         Red_SubCellInst_LFInst_5_LFInst_1_n1,
         Red_SubCellInst_LFInst_5_LFInst_2_n6,
         Red_SubCellInst_LFInst_5_LFInst_2_n5,
         Red_SubCellInst_LFInst_5_LFInst_2_n4,
         Red_SubCellInst_LFInst_5_LFInst_2_n3,
         Red_SubCellInst_LFInst_5_LFInst_2_n2,
         Red_SubCellInst_LFInst_5_LFInst_2_n1,
         Red_SubCellInst_LFInst_6_LFInst_0_n2,
         Red_SubCellInst_LFInst_6_LFInst_0_n1,
         Red_SubCellInst_LFInst_6_LFInst_1_n4,
         Red_SubCellInst_LFInst_6_LFInst_1_n3,
         Red_SubCellInst_LFInst_6_LFInst_1_n2,
         Red_SubCellInst_LFInst_6_LFInst_1_n1,
         Red_SubCellInst_LFInst_6_LFInst_2_n6,
         Red_SubCellInst_LFInst_6_LFInst_2_n5,
         Red_SubCellInst_LFInst_6_LFInst_2_n4,
         Red_SubCellInst_LFInst_6_LFInst_2_n3,
         Red_SubCellInst_LFInst_6_LFInst_2_n2,
         Red_SubCellInst_LFInst_6_LFInst_2_n1,
         Red_SubCellInst_LFInst_7_LFInst_0_n2,
         Red_SubCellInst_LFInst_7_LFInst_0_n1,
         Red_SubCellInst_LFInst_7_LFInst_1_n4,
         Red_SubCellInst_LFInst_7_LFInst_1_n3,
         Red_SubCellInst_LFInst_7_LFInst_1_n2,
         Red_SubCellInst_LFInst_7_LFInst_1_n1,
         Red_SubCellInst_LFInst_7_LFInst_2_n6,
         Red_SubCellInst_LFInst_7_LFInst_2_n5,
         Red_SubCellInst_LFInst_7_LFInst_2_n4,
         Red_SubCellInst_LFInst_7_LFInst_2_n3,
         Red_SubCellInst_LFInst_7_LFInst_2_n2,
         Red_SubCellInst_LFInst_7_LFInst_2_n1,
         Red_SubCellInst_LFInst_8_LFInst_0_n2,
         Red_SubCellInst_LFInst_8_LFInst_0_n1,
         Red_SubCellInst_LFInst_8_LFInst_1_n4,
         Red_SubCellInst_LFInst_8_LFInst_1_n3,
         Red_SubCellInst_LFInst_8_LFInst_1_n2,
         Red_SubCellInst_LFInst_8_LFInst_1_n1,
         Red_SubCellInst_LFInst_8_LFInst_2_n6,
         Red_SubCellInst_LFInst_8_LFInst_2_n5,
         Red_SubCellInst_LFInst_8_LFInst_2_n4,
         Red_SubCellInst_LFInst_8_LFInst_2_n3,
         Red_SubCellInst_LFInst_8_LFInst_2_n2,
         Red_SubCellInst_LFInst_8_LFInst_2_n1,
         Red_SubCellInst_LFInst_9_LFInst_0_n2,
         Red_SubCellInst_LFInst_9_LFInst_0_n1,
         Red_SubCellInst_LFInst_9_LFInst_1_n4,
         Red_SubCellInst_LFInst_9_LFInst_1_n3,
         Red_SubCellInst_LFInst_9_LFInst_1_n2,
         Red_SubCellInst_LFInst_9_LFInst_1_n1,
         Red_SubCellInst_LFInst_9_LFInst_2_n6,
         Red_SubCellInst_LFInst_9_LFInst_2_n5,
         Red_SubCellInst_LFInst_9_LFInst_2_n4,
         Red_SubCellInst_LFInst_9_LFInst_2_n3,
         Red_SubCellInst_LFInst_9_LFInst_2_n2,
         Red_SubCellInst_LFInst_9_LFInst_2_n1,
         Red_SubCellInst_LFInst_10_LFInst_0_n2,
         Red_SubCellInst_LFInst_10_LFInst_0_n1,
         Red_SubCellInst_LFInst_10_LFInst_1_n4,
         Red_SubCellInst_LFInst_10_LFInst_1_n3,
         Red_SubCellInst_LFInst_10_LFInst_1_n2,
         Red_SubCellInst_LFInst_10_LFInst_1_n1,
         Red_SubCellInst_LFInst_10_LFInst_2_n6,
         Red_SubCellInst_LFInst_10_LFInst_2_n5,
         Red_SubCellInst_LFInst_10_LFInst_2_n4,
         Red_SubCellInst_LFInst_10_LFInst_2_n3,
         Red_SubCellInst_LFInst_10_LFInst_2_n2,
         Red_SubCellInst_LFInst_10_LFInst_2_n1,
         Red_SubCellInst_LFInst_11_LFInst_0_n2,
         Red_SubCellInst_LFInst_11_LFInst_0_n1,
         Red_SubCellInst_LFInst_11_LFInst_1_n4,
         Red_SubCellInst_LFInst_11_LFInst_1_n3,
         Red_SubCellInst_LFInst_11_LFInst_1_n2,
         Red_SubCellInst_LFInst_11_LFInst_1_n1,
         Red_SubCellInst_LFInst_11_LFInst_2_n6,
         Red_SubCellInst_LFInst_11_LFInst_2_n5,
         Red_SubCellInst_LFInst_11_LFInst_2_n4,
         Red_SubCellInst_LFInst_11_LFInst_2_n3,
         Red_SubCellInst_LFInst_11_LFInst_2_n2,
         Red_SubCellInst_LFInst_11_LFInst_2_n1,
         Red_SubCellInst_LFInst_12_LFInst_0_n2,
         Red_SubCellInst_LFInst_12_LFInst_0_n1,
         Red_SubCellInst_LFInst_12_LFInst_1_n4,
         Red_SubCellInst_LFInst_12_LFInst_1_n3,
         Red_SubCellInst_LFInst_12_LFInst_1_n2,
         Red_SubCellInst_LFInst_12_LFInst_1_n1,
         Red_SubCellInst_LFInst_12_LFInst_2_n6,
         Red_SubCellInst_LFInst_12_LFInst_2_n5,
         Red_SubCellInst_LFInst_12_LFInst_2_n4,
         Red_SubCellInst_LFInst_12_LFInst_2_n3,
         Red_SubCellInst_LFInst_12_LFInst_2_n2,
         Red_SubCellInst_LFInst_12_LFInst_2_n1,
         Red_SubCellInst_LFInst_13_LFInst_0_n2,
         Red_SubCellInst_LFInst_13_LFInst_0_n1,
         Red_SubCellInst_LFInst_13_LFInst_1_n4,
         Red_SubCellInst_LFInst_13_LFInst_1_n3,
         Red_SubCellInst_LFInst_13_LFInst_1_n2,
         Red_SubCellInst_LFInst_13_LFInst_1_n1,
         Red_SubCellInst_LFInst_13_LFInst_2_n6,
         Red_SubCellInst_LFInst_13_LFInst_2_n5,
         Red_SubCellInst_LFInst_13_LFInst_2_n4,
         Red_SubCellInst_LFInst_13_LFInst_2_n3,
         Red_SubCellInst_LFInst_13_LFInst_2_n2,
         Red_SubCellInst_LFInst_13_LFInst_2_n1,
         Red_SubCellInst_LFInst_14_LFInst_0_n2,
         Red_SubCellInst_LFInst_14_LFInst_0_n1,
         Red_SubCellInst_LFInst_14_LFInst_1_n4,
         Red_SubCellInst_LFInst_14_LFInst_1_n3,
         Red_SubCellInst_LFInst_14_LFInst_1_n2,
         Red_SubCellInst_LFInst_14_LFInst_1_n1,
         Red_SubCellInst_LFInst_14_LFInst_2_n6,
         Red_SubCellInst_LFInst_14_LFInst_2_n5,
         Red_SubCellInst_LFInst_14_LFInst_2_n4,
         Red_SubCellInst_LFInst_14_LFInst_2_n3,
         Red_SubCellInst_LFInst_14_LFInst_2_n2,
         Red_SubCellInst_LFInst_14_LFInst_2_n1,
         Red_SubCellInst_LFInst_15_LFInst_0_n2,
         Red_SubCellInst_LFInst_15_LFInst_0_n1,
         Red_SubCellInst_LFInst_15_LFInst_1_n4,
         Red_SubCellInst_LFInst_15_LFInst_1_n3,
         Red_SubCellInst_LFInst_15_LFInst_1_n2,
         Red_SubCellInst_LFInst_15_LFInst_1_n1,
         Red_SubCellInst_LFInst_15_LFInst_2_n6,
         Red_SubCellInst_LFInst_15_LFInst_2_n5,
         Red_SubCellInst_LFInst_15_LFInst_2_n4,
         Red_SubCellInst_LFInst_15_LFInst_2_n3,
         Red_SubCellInst_LFInst_15_LFInst_2_n2,
         Red_SubCellInst_LFInst_15_LFInst_2_n1, KeyMUX_n3, KeyMUX_n2,
         KeyMUX_n1, Red_K0Inst_LFInst_0_LFInst_0_n1,
         Red_K0Inst_LFInst_0_LFInst_1_n1, Red_K0Inst_LFInst_0_LFInst_2_n1,
         Red_K0Inst_LFInst_1_LFInst_0_n1, Red_K0Inst_LFInst_1_LFInst_1_n1,
         Red_K0Inst_LFInst_1_LFInst_2_n1, Red_K0Inst_LFInst_2_LFInst_0_n1,
         Red_K0Inst_LFInst_2_LFInst_1_n1, Red_K0Inst_LFInst_2_LFInst_2_n1,
         Red_K0Inst_LFInst_3_LFInst_0_n1, Red_K0Inst_LFInst_3_LFInst_1_n1,
         Red_K0Inst_LFInst_3_LFInst_2_n1, Red_K0Inst_LFInst_4_LFInst_0_n1,
         Red_K0Inst_LFInst_4_LFInst_1_n1, Red_K0Inst_LFInst_4_LFInst_2_n1,
         Red_K0Inst_LFInst_5_LFInst_0_n1, Red_K0Inst_LFInst_5_LFInst_1_n1,
         Red_K0Inst_LFInst_5_LFInst_2_n1, Red_K0Inst_LFInst_6_LFInst_0_n1,
         Red_K0Inst_LFInst_6_LFInst_1_n1, Red_K0Inst_LFInst_6_LFInst_2_n1,
         Red_K0Inst_LFInst_7_LFInst_0_n1, Red_K0Inst_LFInst_7_LFInst_1_n1,
         Red_K0Inst_LFInst_7_LFInst_2_n1, Red_K0Inst_LFInst_8_LFInst_0_n1,
         Red_K0Inst_LFInst_8_LFInst_1_n1, Red_K0Inst_LFInst_8_LFInst_2_n1,
         Red_K0Inst_LFInst_9_LFInst_0_n1, Red_K0Inst_LFInst_9_LFInst_1_n1,
         Red_K0Inst_LFInst_9_LFInst_2_n1, Red_K0Inst_LFInst_10_LFInst_0_n1,
         Red_K0Inst_LFInst_10_LFInst_1_n1, Red_K0Inst_LFInst_10_LFInst_2_n1,
         Red_K0Inst_LFInst_11_LFInst_0_n1, Red_K0Inst_LFInst_11_LFInst_1_n1,
         Red_K0Inst_LFInst_11_LFInst_2_n1, Red_K0Inst_LFInst_12_LFInst_0_n1,
         Red_K0Inst_LFInst_12_LFInst_1_n1, Red_K0Inst_LFInst_12_LFInst_2_n1,
         Red_K0Inst_LFInst_13_LFInst_0_n1, Red_K0Inst_LFInst_13_LFInst_1_n1,
         Red_K0Inst_LFInst_13_LFInst_2_n1, Red_K0Inst_LFInst_14_LFInst_0_n1,
         Red_K0Inst_LFInst_14_LFInst_1_n1, Red_K0Inst_LFInst_14_LFInst_2_n1,
         Red_K0Inst_LFInst_15_LFInst_0_n1, Red_K0Inst_LFInst_15_LFInst_1_n1,
         Red_K0Inst_LFInst_15_LFInst_2_n1, Red_K1Inst_LFInst_0_LFInst_0_n1,
         Red_K1Inst_LFInst_0_LFInst_1_n1, Red_K1Inst_LFInst_0_LFInst_2_n1,
         Red_K1Inst_LFInst_1_LFInst_0_n1, Red_K1Inst_LFInst_1_LFInst_1_n1,
         Red_K1Inst_LFInst_1_LFInst_2_n1, Red_K1Inst_LFInst_2_LFInst_0_n1,
         Red_K1Inst_LFInst_2_LFInst_1_n1, Red_K1Inst_LFInst_2_LFInst_2_n1,
         Red_K1Inst_LFInst_3_LFInst_0_n1, Red_K1Inst_LFInst_3_LFInst_1_n1,
         Red_K1Inst_LFInst_3_LFInst_2_n1, Red_K1Inst_LFInst_4_LFInst_0_n1,
         Red_K1Inst_LFInst_4_LFInst_1_n1, Red_K1Inst_LFInst_4_LFInst_2_n1,
         Red_K1Inst_LFInst_5_LFInst_0_n1, Red_K1Inst_LFInst_5_LFInst_1_n1,
         Red_K1Inst_LFInst_5_LFInst_2_n1, Red_K1Inst_LFInst_6_LFInst_0_n1,
         Red_K1Inst_LFInst_6_LFInst_1_n1, Red_K1Inst_LFInst_6_LFInst_2_n1,
         Red_K1Inst_LFInst_7_LFInst_0_n1, Red_K1Inst_LFInst_7_LFInst_1_n1,
         Red_K1Inst_LFInst_7_LFInst_2_n1, Red_K1Inst_LFInst_8_LFInst_0_n1,
         Red_K1Inst_LFInst_8_LFInst_1_n1, Red_K1Inst_LFInst_8_LFInst_2_n1,
         Red_K1Inst_LFInst_9_LFInst_0_n1, Red_K1Inst_LFInst_9_LFInst_1_n1,
         Red_K1Inst_LFInst_9_LFInst_2_n1, Red_K1Inst_LFInst_10_LFInst_0_n1,
         Red_K1Inst_LFInst_10_LFInst_1_n1, Red_K1Inst_LFInst_10_LFInst_2_n1,
         Red_K1Inst_LFInst_11_LFInst_0_n1, Red_K1Inst_LFInst_11_LFInst_1_n1,
         Red_K1Inst_LFInst_11_LFInst_2_n1, Red_K1Inst_LFInst_12_LFInst_0_n1,
         Red_K1Inst_LFInst_12_LFInst_1_n1, Red_K1Inst_LFInst_12_LFInst_2_n1,
         Red_K1Inst_LFInst_13_LFInst_0_n1, Red_K1Inst_LFInst_13_LFInst_1_n1,
         Red_K1Inst_LFInst_13_LFInst_2_n1, Red_K1Inst_LFInst_14_LFInst_0_n1,
         Red_K1Inst_LFInst_14_LFInst_1_n1, Red_K1Inst_LFInst_14_LFInst_2_n1,
         Red_K1Inst_LFInst_15_LFInst_0_n1, Red_K1Inst_LFInst_15_LFInst_1_n1,
         Red_K1Inst_LFInst_15_LFInst_2_n1, Red_KeyMUX_n6, Red_KeyMUX_n5,
         Red_KeyMUX_n4, Red_KeyMUX_n3, Red_KeyMUX_n2, Red_KeyMUX_n1,
         Red_KeyMUX_MUX2to1Inst_0_S_2__0_, Red_KeyMUX_MUX2to1Inst_0_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_0_S_1__0_, Red_KeyMUX_MUX2to1Inst_1_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_1_S_1__1_, Red_KeyMUX_MUX2to1Inst_1_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_2_S_2__0_, Red_KeyMUX_MUX2to1Inst_2_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_2_S_1__0_, Red_KeyMUX_MUX2to1Inst_3_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_3_S_1__1_, Red_KeyMUX_MUX2to1Inst_3_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_4_S_2__0_, Red_KeyMUX_MUX2to1Inst_4_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_4_S_1__0_, Red_KeyMUX_MUX2to1Inst_5_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_5_S_1__1_, Red_KeyMUX_MUX2to1Inst_5_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_6_S_2__0_, Red_KeyMUX_MUX2to1Inst_6_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_6_S_1__0_, Red_KeyMUX_MUX2to1Inst_7_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_7_S_1__1_, Red_KeyMUX_MUX2to1Inst_7_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_8_S_2__0_, Red_KeyMUX_MUX2to1Inst_8_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_8_S_1__0_, Red_KeyMUX_MUX2to1Inst_9_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_9_S_1__1_, Red_KeyMUX_MUX2to1Inst_9_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_10_S_2__0_, Red_KeyMUX_MUX2to1Inst_10_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_10_S_1__0_, Red_KeyMUX_MUX2to1Inst_11_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_11_S_1__1_, Red_KeyMUX_MUX2to1Inst_11_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_12_S_2__0_, Red_KeyMUX_MUX2to1Inst_12_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_12_S_1__0_, Red_KeyMUX_MUX2to1Inst_13_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_13_S_1__1_, Red_KeyMUX_MUX2to1Inst_13_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_14_S_2__0_, Red_KeyMUX_MUX2to1Inst_14_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_14_S_1__0_, Red_KeyMUX_MUX2to1Inst_15_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_15_S_1__1_, Red_KeyMUX_MUX2to1Inst_15_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_16_S_2__0_, Red_KeyMUX_MUX2to1Inst_16_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_16_S_1__0_, Red_KeyMUX_MUX2to1Inst_17_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_17_S_1__1_, Red_KeyMUX_MUX2to1Inst_17_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_18_S_2__0_, Red_KeyMUX_MUX2to1Inst_18_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_18_S_1__0_, Red_KeyMUX_MUX2to1Inst_19_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_19_S_1__1_, Red_KeyMUX_MUX2to1Inst_19_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_20_S_2__0_, Red_KeyMUX_MUX2to1Inst_20_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_20_S_1__0_, Red_KeyMUX_MUX2to1Inst_21_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_21_S_1__1_, Red_KeyMUX_MUX2to1Inst_21_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_22_S_2__0_, Red_KeyMUX_MUX2to1Inst_22_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_22_S_1__0_, Red_KeyMUX_MUX2to1Inst_23_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_23_S_1__1_, Red_KeyMUX_MUX2to1Inst_23_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_24_S_2__0_, Red_KeyMUX_MUX2to1Inst_24_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_24_S_1__0_, Red_KeyMUX_MUX2to1Inst_25_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_25_S_1__1_, Red_KeyMUX_MUX2to1Inst_25_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_26_S_2__0_, Red_KeyMUX_MUX2to1Inst_26_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_26_S_1__0_, Red_KeyMUX_MUX2to1Inst_27_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_27_S_1__1_, Red_KeyMUX_MUX2to1Inst_27_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_28_S_2__0_, Red_KeyMUX_MUX2to1Inst_28_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_28_S_1__0_, Red_KeyMUX_MUX2to1Inst_29_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_29_S_1__1_, Red_KeyMUX_MUX2to1Inst_29_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_30_S_2__0_, Red_KeyMUX_MUX2to1Inst_30_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_30_S_1__0_, Red_KeyMUX_MUX2to1Inst_31_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_31_S_1__1_, Red_KeyMUX_MUX2to1Inst_31_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_32_S_2__0_, Red_KeyMUX_MUX2to1Inst_32_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_32_S_1__0_, Red_KeyMUX_MUX2to1Inst_33_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_33_S_1__1_, Red_KeyMUX_MUX2to1Inst_33_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_34_S_2__0_, Red_KeyMUX_MUX2to1Inst_34_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_34_S_1__0_, Red_KeyMUX_MUX2to1Inst_35_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_35_S_1__1_, Red_KeyMUX_MUX2to1Inst_35_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_36_S_2__0_, Red_KeyMUX_MUX2to1Inst_36_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_36_S_1__0_, Red_KeyMUX_MUX2to1Inst_37_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_37_S_1__1_, Red_KeyMUX_MUX2to1Inst_37_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_38_S_2__0_, Red_KeyMUX_MUX2to1Inst_38_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_38_S_1__0_, Red_KeyMUX_MUX2to1Inst_39_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_39_S_1__1_, Red_KeyMUX_MUX2to1Inst_39_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_40_S_2__0_, Red_KeyMUX_MUX2to1Inst_40_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_40_S_1__0_, Red_KeyMUX_MUX2to1Inst_41_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_41_S_1__1_, Red_KeyMUX_MUX2to1Inst_41_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_42_S_2__0_, Red_KeyMUX_MUX2to1Inst_42_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_42_S_1__0_, Red_KeyMUX_MUX2to1Inst_43_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_43_S_1__1_, Red_KeyMUX_MUX2to1Inst_43_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_44_S_2__0_, Red_KeyMUX_MUX2to1Inst_44_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_44_S_1__0_, Red_KeyMUX_MUX2to1Inst_45_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_45_S_1__1_, Red_KeyMUX_MUX2to1Inst_45_S_1__0_,
         Red_KeyMUX_MUX2to1Inst_46_S_2__0_, Red_KeyMUX_MUX2to1Inst_46_S_1__1_,
         Red_KeyMUX_MUX2to1Inst_46_S_1__0_, Red_KeyMUX_MUX2to1Inst_47_S_2__0_,
         Red_KeyMUX_MUX2to1Inst_47_S_1__1_, Red_KeyMUX_MUX2to1Inst_47_S_1__0_,
         FSMSignals_doneInst_n1, Red_FSMUpdateInst_Red_StateUpdateBitInst_2_n1,
         Red_FSMUpdateInst_Red_StateUpdateBitInst_3_n1,
         Red_FSMUpdateInst_Red_StateUpdateBitInst_5_n2,
         Red_FSMUpdateInst_Red_StateUpdateBitInst_5_n1,
         Red_FSMSignals_doneInst_Red_FSMSignals_doneBitInst_0_n1,
         Red_FSMSignals_doneInst_Red_FSMSignals_doneBitInst_1_n1,
         Red_ToCheckInst_LFInst_0_LFInst_0_n1,
         Red_ToCheckInst_LFInst_0_LFInst_1_n1,
         Red_ToCheckInst_LFInst_0_LFInst_2_n1,
         Red_ToCheckInst_LFInst_1_LFInst_0_n1,
         Red_ToCheckInst_LFInst_1_LFInst_1_n1,
         Red_ToCheckInst_LFInst_1_LFInst_2_n1,
         Red_ToCheckInst_LFInst_2_LFInst_0_n1,
         Red_ToCheckInst_LFInst_2_LFInst_1_n1,
         Red_ToCheckInst_LFInst_2_LFInst_2_n1,
         Red_ToCheckInst_LFInst_3_LFInst_0_n1,
         Red_ToCheckInst_LFInst_3_LFInst_1_n1,
         Red_ToCheckInst_LFInst_3_LFInst_2_n1,
         Red_ToCheckInst_LFInst_4_LFInst_0_n1,
         Red_ToCheckInst_LFInst_4_LFInst_1_n1,
         Red_ToCheckInst_LFInst_4_LFInst_2_n1,
         Red_ToCheckInst_LFInst_5_LFInst_0_n1,
         Red_ToCheckInst_LFInst_5_LFInst_1_n1,
         Red_ToCheckInst_LFInst_5_LFInst_2_n1,
         Red_ToCheckInst_LFInst_6_LFInst_0_n1,
         Red_ToCheckInst_LFInst_6_LFInst_1_n1,
         Red_ToCheckInst_LFInst_6_LFInst_2_n1,
         Red_ToCheckInst_LFInst_7_LFInst_0_n1,
         Red_ToCheckInst_LFInst_7_LFInst_1_n1,
         Red_ToCheckInst_LFInst_7_LFInst_2_n1,
         Red_ToCheckInst_LFInst_8_LFInst_0_n1,
         Red_ToCheckInst_LFInst_8_LFInst_1_n1,
         Red_ToCheckInst_LFInst_8_LFInst_2_n1,
         Red_ToCheckInst_LFInst_9_LFInst_0_n1,
         Red_ToCheckInst_LFInst_9_LFInst_1_n1,
         Red_ToCheckInst_LFInst_9_LFInst_2_n1,
         Red_ToCheckInst_LFInst_10_LFInst_0_n1,
         Red_ToCheckInst_LFInst_10_LFInst_1_n1,
         Red_ToCheckInst_LFInst_10_LFInst_2_n1,
         Red_ToCheckInst_LFInst_11_LFInst_0_n1,
         Red_ToCheckInst_LFInst_11_LFInst_1_n1,
         Red_ToCheckInst_LFInst_11_LFInst_2_n1,
         Red_ToCheckInst_LFInst_12_LFInst_0_n1,
         Red_ToCheckInst_LFInst_12_LFInst_1_n1,
         Red_ToCheckInst_LFInst_12_LFInst_2_n1,
         Red_ToCheckInst_LFInst_13_LFInst_0_n1,
         Red_ToCheckInst_LFInst_13_LFInst_1_n1,
         Red_ToCheckInst_LFInst_13_LFInst_2_n1,
         Red_ToCheckInst_LFInst_14_LFInst_0_n1,
         Red_ToCheckInst_LFInst_14_LFInst_1_n1,
         Red_ToCheckInst_LFInst_14_LFInst_2_n1,
         Red_ToCheckInst_LFInst_15_LFInst_0_n1,
         Red_ToCheckInst_LFInst_15_LFInst_1_n1,
         Red_ToCheckInst_LFInst_15_LFInst_2_n1,
         Red_ToCheckInst_LFInst_16_LFInst_0_n1,
         Red_ToCheckInst_LFInst_16_LFInst_1_n1,
         Red_ToCheckInst_LFInst_16_LFInst_2_n1,
         Red_ToCheckInst_LFInst_17_LFInst_0_n1,
         Red_ToCheckInst_LFInst_17_LFInst_1_n1,
         Red_ToCheckInst_LFInst_17_LFInst_2_n1,
         Red_ToCheckInst_LFInst_18_LFInst_0_n1,
         Red_ToCheckInst_LFInst_18_LFInst_1_n1,
         Red_ToCheckInst_LFInst_18_LFInst_2_n1,
         Red_ToCheckInst_LFInst_19_LFInst_0_n1,
         Red_ToCheckInst_LFInst_19_LFInst_1_n1,
         Red_ToCheckInst_LFInst_19_LFInst_2_n1,
         Red_ToCheckInst_LFInst_20_LFInst_0_n1,
         Red_ToCheckInst_LFInst_20_LFInst_1_n1,
         Red_ToCheckInst_LFInst_20_LFInst_2_n1,
         Red_ToCheckInst_LFInst_21_LFInst_0_n1,
         Red_ToCheckInst_LFInst_21_LFInst_1_n1,
         Red_ToCheckInst_LFInst_21_LFInst_2_n1,
         Red_ToCheckInst_LFInst_22_LFInst_0_n1,
         Red_ToCheckInst_LFInst_22_LFInst_1_n1,
         Red_ToCheckInst_LFInst_22_LFInst_2_n1,
         Red_ToCheckInst_LFInst_23_LFInst_0_n1,
         Red_ToCheckInst_LFInst_23_LFInst_1_n1,
         Red_ToCheckInst_LFInst_23_LFInst_2_n1,
         Red_ToCheckInst_LFInst_24_LFInst_0_n1,
         Red_ToCheckInst_LFInst_24_LFInst_1_n1,
         Red_ToCheckInst_LFInst_24_LFInst_2_n1,
         Red_ToCheckInst_LFInst_25_LFInst_0_n1,
         Red_ToCheckInst_LFInst_25_LFInst_1_n1,
         Red_ToCheckInst_LFInst_25_LFInst_2_n1,
         Red_ToCheckInst_LFInst_26_LFInst_0_n1,
         Red_ToCheckInst_LFInst_26_LFInst_1_n1,
         Red_ToCheckInst_LFInst_26_LFInst_2_n1,
         Red_ToCheckInst_LFInst_27_LFInst_0_n1,
         Red_ToCheckInst_LFInst_27_LFInst_1_n1,
         Red_ToCheckInst_LFInst_27_LFInst_2_n1,
         Red_ToCheckInst_LFInst_28_LFInst_0_n1,
         Red_ToCheckInst_LFInst_28_LFInst_1_n1,
         Red_ToCheckInst_LFInst_28_LFInst_2_n1,
         Red_ToCheckInst_LFInst_29_LFInst_0_n1,
         Red_ToCheckInst_LFInst_29_LFInst_1_n1,
         Red_ToCheckInst_LFInst_29_LFInst_2_n1,
         Red_ToCheckInst_LFInst_30_LFInst_0_n1,
         Red_ToCheckInst_LFInst_30_LFInst_1_n1,
         Red_ToCheckInst_LFInst_30_LFInst_2_n1,
         Red_ToCheckInst_LFInst_31_LFInst_0_n1,
         Red_ToCheckInst_LFInst_31_LFInst_1_n1,
         Red_ToCheckInst_LFInst_31_LFInst_2_n1,
         Red_ToCheckInst_LFInst_32_LFInst_0_n1,
         Red_ToCheckInst_LFInst_32_LFInst_1_n1,
         Red_ToCheckInst_LFInst_32_LFInst_2_n1,
         Red_ToCheckInst_LFInst_33_LFInst_0_n1,
         Red_ToCheckInst_LFInst_33_LFInst_1_n1,
         Red_ToCheckInst_LFInst_33_LFInst_2_n1,
         Red_ToCheckInst_LFInst_34_LFInst_0_n1,
         Red_ToCheckInst_LFInst_34_LFInst_1_n1,
         Red_ToCheckInst_LFInst_34_LFInst_2_n1,
         Red_ToCheckInst_LFInst_35_LFInst_0_n1,
         Red_ToCheckInst_LFInst_35_LFInst_1_n1,
         Red_ToCheckInst_LFInst_35_LFInst_2_n1,
         Red_ToCheckInst_LFInst_36_LFInst_0_n1,
         Red_ToCheckInst_LFInst_36_LFInst_1_n1,
         Red_ToCheckInst_LFInst_36_LFInst_2_n1,
         Red_ToCheckInst_LFInst_37_LFInst_0_n1,
         Red_ToCheckInst_LFInst_37_LFInst_1_n1,
         Red_ToCheckInst_LFInst_37_LFInst_2_n1,
         Red_ToCheckInst_LFInst_38_LFInst_0_n1,
         Red_ToCheckInst_LFInst_38_LFInst_1_n1,
         Red_ToCheckInst_LFInst_38_LFInst_2_n1,
         Red_ToCheckInst_LFInst_39_LFInst_0_n1,
         Red_ToCheckInst_LFInst_39_LFInst_1_n1,
         Red_ToCheckInst_LFInst_39_LFInst_2_n1,
         Red_ToCheckInst_LFInst_40_LFInst_0_n1,
         Red_ToCheckInst_LFInst_40_LFInst_1_n1,
         Red_ToCheckInst_LFInst_40_LFInst_2_n1, Check1_CheckInst_0_n54,
         Check1_CheckInst_0_n53, Check1_CheckInst_0_n52,
         Check1_CheckInst_0_n51, Check1_CheckInst_0_n50,
         Check1_CheckInst_0_n49, Check1_CheckInst_0_n48,
         Check1_CheckInst_0_n47, Check1_CheckInst_0_n46,
         Check1_CheckInst_0_n45, Check1_CheckInst_0_n44,
         Check1_CheckInst_0_n43, Check1_CheckInst_0_n42,
         Check1_CheckInst_0_n41, Check1_CheckInst_0_n40,
         Check1_CheckInst_0_n39, Check1_CheckInst_0_n38,
         Check1_CheckInst_0_n37, Check1_CheckInst_0_n36,
         Check1_CheckInst_0_n35, Check1_CheckInst_0_n34,
         Check1_CheckInst_0_n33, Check1_CheckInst_0_n32,
         Check1_CheckInst_0_n31, Check1_CheckInst_0_n30,
         Check1_CheckInst_0_n29, Check1_CheckInst_0_n28,
         Check1_CheckInst_0_n27, Check1_CheckInst_0_n26,
         Check1_CheckInst_0_n25, Check1_CheckInst_0_n24,
         Check1_CheckInst_0_n23, Check1_CheckInst_0_n22,
         Check1_CheckInst_0_n21, Check1_CheckInst_0_n20,
         Check1_CheckInst_0_n19, Check1_CheckInst_0_n18,
         Check1_CheckInst_0_n17, Check1_CheckInst_0_n16,
         Check1_CheckInst_0_n15, Check1_CheckInst_0_n14,
         Check1_CheckInst_0_n13, Check1_CheckInst_0_n12,
         Check1_CheckInst_0_n11, Check1_CheckInst_0_n10, Check1_CheckInst_0_n9,
         Check1_CheckInst_0_n8, Check1_CheckInst_0_n7, Check1_CheckInst_0_n6,
         Check1_CheckInst_0_n5, Check1_CheckInst_0_n4, Check1_CheckInst_0_n3,
         Check1_CheckInst_0_n2, Check1_CheckInst_0_n1, Check1_CheckInst_1_n54,
         Check1_CheckInst_1_n53, Check1_CheckInst_1_n52,
         Check1_CheckInst_1_n51, Check1_CheckInst_1_n50,
         Check1_CheckInst_1_n49, Check1_CheckInst_1_n48,
         Check1_CheckInst_1_n47, Check1_CheckInst_1_n46,
         Check1_CheckInst_1_n45, Check1_CheckInst_1_n44,
         Check1_CheckInst_1_n43, Check1_CheckInst_1_n42,
         Check1_CheckInst_1_n41, Check1_CheckInst_1_n40,
         Check1_CheckInst_1_n39, Check1_CheckInst_1_n38,
         Check1_CheckInst_1_n37, Check1_CheckInst_1_n36,
         Check1_CheckInst_1_n35, Check1_CheckInst_1_n34,
         Check1_CheckInst_1_n33, Check1_CheckInst_1_n32,
         Check1_CheckInst_1_n31, Check1_CheckInst_1_n30,
         Check1_CheckInst_1_n29, Check1_CheckInst_1_n28,
         Check1_CheckInst_1_n27, Check1_CheckInst_1_n26,
         Check1_CheckInst_1_n25, Check1_CheckInst_1_n24,
         Check1_CheckInst_1_n23, Check1_CheckInst_1_n22,
         Check1_CheckInst_1_n21, Check1_CheckInst_1_n20,
         Check1_CheckInst_1_n19, Check1_CheckInst_1_n18,
         Check1_CheckInst_1_n17, Check1_CheckInst_1_n16,
         Check1_CheckInst_1_n15, Check1_CheckInst_1_n14,
         Check1_CheckInst_1_n13, Check1_CheckInst_1_n12,
         Check1_CheckInst_1_n11, Check1_CheckInst_1_n10, Check1_CheckInst_1_n9,
         Check1_CheckInst_1_n8, Check1_CheckInst_1_n7, Check1_CheckInst_1_n6,
         Check1_CheckInst_1_n5, Check1_CheckInst_1_n4, Check1_CheckInst_1_n3,
         Check1_CheckInst_1_n2, Check1_CheckInst_1_n1, Check1_CheckInst_2_n54,
         Check1_CheckInst_2_n53, Check1_CheckInst_2_n52,
         Check1_CheckInst_2_n51, Check1_CheckInst_2_n50,
         Check1_CheckInst_2_n49, Check1_CheckInst_2_n48,
         Check1_CheckInst_2_n47, Check1_CheckInst_2_n46,
         Check1_CheckInst_2_n45, Check1_CheckInst_2_n44,
         Check1_CheckInst_2_n43, Check1_CheckInst_2_n42,
         Check1_CheckInst_2_n41, Check1_CheckInst_2_n40,
         Check1_CheckInst_2_n39, Check1_CheckInst_2_n38,
         Check1_CheckInst_2_n37, Check1_CheckInst_2_n36,
         Check1_CheckInst_2_n35, Check1_CheckInst_2_n34,
         Check1_CheckInst_2_n33, Check1_CheckInst_2_n32,
         Check1_CheckInst_2_n31, Check1_CheckInst_2_n30,
         Check1_CheckInst_2_n29, Check1_CheckInst_2_n28,
         Check1_CheckInst_2_n27, Check1_CheckInst_2_n26,
         Check1_CheckInst_2_n25, Check1_CheckInst_2_n24,
         Check1_CheckInst_2_n23, Check1_CheckInst_2_n22,
         Check1_CheckInst_2_n21, Check1_CheckInst_2_n20,
         Check1_CheckInst_2_n19, Check1_CheckInst_2_n18,
         Check1_CheckInst_2_n17, Check1_CheckInst_2_n16,
         Check1_CheckInst_2_n15, Check1_CheckInst_2_n14,
         Check1_CheckInst_2_n13, Check1_CheckInst_2_n12,
         Check1_CheckInst_2_n11, Check1_CheckInst_2_n10, Check1_CheckInst_2_n9,
         Check1_CheckInst_2_n8, Check1_CheckInst_2_n7, Check1_CheckInst_2_n6,
         Check1_CheckInst_2_n5, Check1_CheckInst_2_n4, Check1_CheckInst_2_n3,
         Check1_CheckInst_2_n2, Check1_CheckInst_2_n1, ANDInst_0_n2,
         ANDInst_0_n1, ANDInst_1_n2, ANDInst_1_n1, ANDInst_2_n2, ANDInst_2_n1,
         ANDInst_3_n2, ANDInst_3_n1, ANDInst_4_n2, ANDInst_4_n1, OutputMUX_n15,
         OutputMUX_n14, OutputMUX_n13, OutputMUX_n12, OutputMUX_n11,
         OutputMUX_n10, OutputMUX_n9, OutputMUX_n8, OutputMUX_n7, OutputMUX_n6,
         OutputMUX_n5, OutputMUX_n4, OutputMUX_n3, OutputMUX_n2, OutputMUX_n1,
         OutputReg_n71, OutputReg_n70, OutputReg_n69, OutputReg_n68,
         OutputReg_n67, OutputReg_n3, OutputReg_n2, OutputReg_n66,
         OutputReg_n65, OutputReg_n64, OutputReg_n63, OutputReg_n62,
         OutputReg_n61, OutputReg_n60, OutputReg_n59, OutputReg_n58,
         OutputReg_n57, OutputReg_n56, OutputReg_n55, OutputReg_n54,
         OutputReg_n53, OutputReg_n52, OutputReg_n51, OutputReg_n50,
         OutputReg_n49, OutputReg_n48, OutputReg_n47, OutputReg_n46,
         OutputReg_n45, OutputReg_n44, OutputReg_n43, OutputReg_n42,
         OutputReg_n41, OutputReg_n40, OutputReg_n39, OutputReg_n38,
         OutputReg_n37, OutputReg_n36, OutputReg_n35, OutputReg_n34,
         OutputReg_n33, OutputReg_n32, OutputReg_n31, OutputReg_n30,
         OutputReg_n29, OutputReg_n28, OutputReg_n27, OutputReg_n26,
         OutputReg_n25, OutputReg_n24, OutputReg_n23, OutputReg_n22,
         OutputReg_n21, OutputReg_n20, OutputReg_n19, OutputReg_n18,
         OutputReg_n17, OutputReg_n16, OutputReg_n15, OutputReg_n14,
         OutputReg_n13, OutputReg_n12, OutputReg_n11, OutputReg_n10,
         OutputReg_n9, OutputReg_n8, OutputReg_n7, OutputReg_n6, OutputReg_n5,
         OutputReg_n4, OutputReg_n1;
  wire   [63:0] Feedback;
  wire   [63:32] MCInput;
  wire   [63:0] MCOutput;
  wire   [63:0] AddRoundKeyOutput;
  wire   [63:0] PermutationOutput;
  wire   [47:0] Red_Input;
  wire   [47:0] Red_Feedback;
  wire   [47:24] Red_MCInput;
  wire   [47:0] Red_MCOutput;
  wire   [5:0] Red_RoundConstant;
  wire   [47:0] Red_StateRegOutput;
  wire   [63:0] SelectedKey;
  wire   [47:0] Red_K0;
  wire   [47:0] Red_K1;
  wire   [2:0] Red_sel_Key;
  wire   [47:0] Red_SelectedKey;
  wire   [6:0] FSMReg;
  wire   [6:0] FSMUpdate;
  wire   [1:0] selects;
  wire   [1:0] selectsReg;
  wire   [1:0] selectsNext;
  wire   [5:0] Red_FSMReg;
  wire   [5:0] Red_FSMUpdate;
  wire   [1:0] Red_done;
  wire   [2:0] Red_sel_Tweak;
  wire   [5:0] Red_selectsReg;
  wire   [4:0] Red_selectsNext;
  wire   [47:0] Red_final;
  wire   [122:0] Red_SignaltoCheck;
  wire   [2:0] Error;
  wire   [4:0] ErrorFree;
  wire   [4:0] ErrorFreeUpdate;
  wire   [63:0] OutputRegIn;
  wire   [4:1] OutputMUX_MUX2to1Inst_0_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_1_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_2_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_3_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_4_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_5_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_6_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_7_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_8_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_9_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_10_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_11_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_12_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_13_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_14_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_15_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_16_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_17_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_18_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_19_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_20_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_21_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_22_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_23_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_24_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_25_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_26_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_27_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_28_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_29_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_30_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_31_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_32_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_33_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_34_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_35_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_36_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_37_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_38_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_39_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_40_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_41_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_42_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_43_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_44_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_45_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_46_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_47_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_48_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_49_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_50_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_51_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_52_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_53_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_54_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_55_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_56_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_57_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_58_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_59_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_60_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_61_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_62_sig;
  wire   [4:1] OutputMUX_MUX2to1Inst_63_sig;

  DFF_X1 ErrorFree_reg_0_ ( .D(N3), .CK(clk), .Q(ErrorFree[0]), .QN() );
  DFF_X1 ErrorFree_reg_1_ ( .D(N4), .CK(clk), .Q(ErrorFree[1]), .QN() );
  DFF_X1 ErrorFree_reg_2_ ( .D(N5), .CK(clk), .Q(ErrorFree[2]), .QN() );
  DFF_X1 ErrorFree_reg_3_ ( .D(N6), .CK(clk), .Q(ErrorFree[3]), .QN() );
  DFF_X1 ErrorFree_reg_4_ ( .D(N7), .CK(clk), .Q(ErrorFree[4]), .QN() );
  OR2_X1 U9 ( .A1(rst), .A2(ErrorFreeUpdate[0]), .ZN(N3) );
  OR2_X1 U10 ( .A1(rst), .A2(ErrorFreeUpdate[1]), .ZN(N4) );
  OR2_X1 U11 ( .A1(rst), .A2(ErrorFreeUpdate[2]), .ZN(N5) );
  OR2_X1 U12 ( .A1(rst), .A2(ErrorFreeUpdate[3]), .ZN(N6) );
  OR2_X1 U13 ( .A1(rst), .A2(ErrorFreeUpdate[4]), .ZN(N7) );
  MUX2_X1 InputMUX_MUXInst_0_U1 ( .A(Feedback[0]), .B(Input[0]), .S(rst), .Z(
        MCOutput[0]) );
  MUX2_X1 InputMUX_MUXInst_1_U1 ( .A(Feedback[1]), .B(Input[1]), .S(rst), .Z(
        MCOutput[1]) );
  MUX2_X1 InputMUX_MUXInst_2_U1 ( .A(Feedback[2]), .B(Input[2]), .S(rst), .Z(
        MCOutput[2]) );
  MUX2_X1 InputMUX_MUXInst_3_U1 ( .A(Feedback[3]), .B(Input[3]), .S(rst), .Z(
        MCOutput[3]) );
  MUX2_X1 InputMUX_MUXInst_4_U1 ( .A(Feedback[4]), .B(Input[4]), .S(rst), .Z(
        MCOutput[4]) );
  MUX2_X1 InputMUX_MUXInst_5_U1 ( .A(Feedback[5]), .B(Input[5]), .S(rst), .Z(
        MCOutput[5]) );
  MUX2_X1 InputMUX_MUXInst_6_U1 ( .A(Feedback[6]), .B(Input[6]), .S(rst), .Z(
        MCOutput[6]) );
  MUX2_X1 InputMUX_MUXInst_7_U1 ( .A(Feedback[7]), .B(Input[7]), .S(rst), .Z(
        MCOutput[7]) );
  MUX2_X1 InputMUX_MUXInst_8_U1 ( .A(Feedback[8]), .B(Input[8]), .S(rst), .Z(
        MCOutput[8]) );
  MUX2_X1 InputMUX_MUXInst_9_U1 ( .A(Feedback[9]), .B(Input[9]), .S(rst), .Z(
        MCOutput[9]) );
  MUX2_X1 InputMUX_MUXInst_10_U1 ( .A(Feedback[10]), .B(Input[10]), .S(rst), 
        .Z(MCOutput[10]) );
  MUX2_X1 InputMUX_MUXInst_11_U1 ( .A(Feedback[11]), .B(Input[11]), .S(rst), 
        .Z(MCOutput[11]) );
  MUX2_X1 InputMUX_MUXInst_12_U1 ( .A(Feedback[12]), .B(Input[12]), .S(rst), 
        .Z(MCOutput[12]) );
  MUX2_X1 InputMUX_MUXInst_13_U1 ( .A(Feedback[13]), .B(Input[13]), .S(rst), 
        .Z(MCOutput[13]) );
  MUX2_X1 InputMUX_MUXInst_14_U1 ( .A(Feedback[14]), .B(Input[14]), .S(rst), 
        .Z(MCOutput[14]) );
  MUX2_X1 InputMUX_MUXInst_15_U1 ( .A(Feedback[15]), .B(Input[15]), .S(rst), 
        .Z(MCOutput[15]) );
  MUX2_X1 InputMUX_MUXInst_16_U1 ( .A(Feedback[16]), .B(Input[16]), .S(rst), 
        .Z(MCOutput[16]) );
  MUX2_X1 InputMUX_MUXInst_17_U1 ( .A(Feedback[17]), .B(Input[17]), .S(rst), 
        .Z(MCOutput[17]) );
  MUX2_X1 InputMUX_MUXInst_18_U1 ( .A(Feedback[18]), .B(Input[18]), .S(rst), 
        .Z(MCOutput[18]) );
  MUX2_X1 InputMUX_MUXInst_19_U1 ( .A(Feedback[19]), .B(Input[19]), .S(rst), 
        .Z(MCOutput[19]) );
  MUX2_X1 InputMUX_MUXInst_20_U1 ( .A(Feedback[20]), .B(Input[20]), .S(rst), 
        .Z(MCOutput[20]) );
  MUX2_X1 InputMUX_MUXInst_21_U1 ( .A(Feedback[21]), .B(Input[21]), .S(rst), 
        .Z(MCOutput[21]) );
  MUX2_X1 InputMUX_MUXInst_22_U1 ( .A(Feedback[22]), .B(Input[22]), .S(rst), 
        .Z(MCOutput[22]) );
  MUX2_X1 InputMUX_MUXInst_23_U1 ( .A(Feedback[23]), .B(Input[23]), .S(rst), 
        .Z(MCOutput[23]) );
  MUX2_X1 InputMUX_MUXInst_24_U1 ( .A(Feedback[24]), .B(Input[24]), .S(rst), 
        .Z(MCOutput[24]) );
  MUX2_X1 InputMUX_MUXInst_25_U1 ( .A(Feedback[25]), .B(Input[25]), .S(rst), 
        .Z(MCOutput[25]) );
  MUX2_X1 InputMUX_MUXInst_26_U1 ( .A(Feedback[26]), .B(Input[26]), .S(rst), 
        .Z(MCOutput[26]) );
  MUX2_X1 InputMUX_MUXInst_27_U1 ( .A(Feedback[27]), .B(Input[27]), .S(rst), 
        .Z(MCOutput[27]) );
  MUX2_X1 InputMUX_MUXInst_28_U1 ( .A(Feedback[28]), .B(Input[28]), .S(rst), 
        .Z(MCOutput[28]) );
  MUX2_X1 InputMUX_MUXInst_29_U1 ( .A(Feedback[29]), .B(Input[29]), .S(rst), 
        .Z(MCOutput[29]) );
  MUX2_X1 InputMUX_MUXInst_30_U1 ( .A(Feedback[30]), .B(Input[30]), .S(rst), 
        .Z(MCOutput[30]) );
  MUX2_X1 InputMUX_MUXInst_31_U1 ( .A(Feedback[31]), .B(Input[31]), .S(rst), 
        .Z(MCOutput[31]) );
  MUX2_X1 InputMUX_MUXInst_32_U1 ( .A(Feedback[32]), .B(Input[32]), .S(rst), 
        .Z(MCInput[32]) );
  MUX2_X1 InputMUX_MUXInst_33_U1 ( .A(Feedback[33]), .B(Input[33]), .S(rst), 
        .Z(MCInput[33]) );
  MUX2_X1 InputMUX_MUXInst_34_U1 ( .A(Feedback[34]), .B(Input[34]), .S(rst), 
        .Z(MCInput[34]) );
  MUX2_X1 InputMUX_MUXInst_35_U1 ( .A(Feedback[35]), .B(Input[35]), .S(rst), 
        .Z(MCInput[35]) );
  MUX2_X1 InputMUX_MUXInst_36_U1 ( .A(Feedback[36]), .B(Input[36]), .S(rst), 
        .Z(MCInput[36]) );
  MUX2_X1 InputMUX_MUXInst_37_U1 ( .A(Feedback[37]), .B(Input[37]), .S(rst), 
        .Z(MCInput[37]) );
  MUX2_X1 InputMUX_MUXInst_38_U1 ( .A(Feedback[38]), .B(Input[38]), .S(rst), 
        .Z(MCInput[38]) );
  MUX2_X1 InputMUX_MUXInst_39_U1 ( .A(Feedback[39]), .B(Input[39]), .S(rst), 
        .Z(MCInput[39]) );
  MUX2_X1 InputMUX_MUXInst_40_U1 ( .A(Feedback[40]), .B(Input[40]), .S(rst), 
        .Z(MCInput[40]) );
  MUX2_X1 InputMUX_MUXInst_41_U1 ( .A(Feedback[41]), .B(Input[41]), .S(rst), 
        .Z(MCInput[41]) );
  MUX2_X1 InputMUX_MUXInst_42_U1 ( .A(Feedback[42]), .B(Input[42]), .S(rst), 
        .Z(MCInput[42]) );
  MUX2_X1 InputMUX_MUXInst_43_U1 ( .A(Feedback[43]), .B(Input[43]), .S(rst), 
        .Z(MCInput[43]) );
  MUX2_X1 InputMUX_MUXInst_44_U1 ( .A(Feedback[44]), .B(Input[44]), .S(rst), 
        .Z(MCInput[44]) );
  MUX2_X1 InputMUX_MUXInst_45_U1 ( .A(Feedback[45]), .B(Input[45]), .S(rst), 
        .Z(MCInput[45]) );
  MUX2_X1 InputMUX_MUXInst_46_U1 ( .A(Feedback[46]), .B(Input[46]), .S(rst), 
        .Z(MCInput[46]) );
  MUX2_X1 InputMUX_MUXInst_47_U1 ( .A(Feedback[47]), .B(Input[47]), .S(rst), 
        .Z(MCInput[47]) );
  MUX2_X1 InputMUX_MUXInst_48_U1 ( .A(Feedback[48]), .B(Input[48]), .S(rst), 
        .Z(MCInput[48]) );
  MUX2_X1 InputMUX_MUXInst_49_U1 ( .A(Feedback[49]), .B(Input[49]), .S(rst), 
        .Z(MCInput[49]) );
  MUX2_X1 InputMUX_MUXInst_50_U1 ( .A(Feedback[50]), .B(Input[50]), .S(rst), 
        .Z(MCInput[50]) );
  MUX2_X1 InputMUX_MUXInst_51_U1 ( .A(Feedback[51]), .B(Input[51]), .S(rst), 
        .Z(MCInput[51]) );
  MUX2_X1 InputMUX_MUXInst_52_U1 ( .A(Feedback[52]), .B(Input[52]), .S(rst), 
        .Z(MCInput[52]) );
  MUX2_X1 InputMUX_MUXInst_53_U1 ( .A(Feedback[53]), .B(Input[53]), .S(rst), 
        .Z(MCInput[53]) );
  MUX2_X1 InputMUX_MUXInst_54_U1 ( .A(Feedback[54]), .B(Input[54]), .S(rst), 
        .Z(MCInput[54]) );
  MUX2_X1 InputMUX_MUXInst_55_U1 ( .A(Feedback[55]), .B(Input[55]), .S(rst), 
        .Z(MCInput[55]) );
  MUX2_X1 InputMUX_MUXInst_56_U1 ( .A(Feedback[56]), .B(Input[56]), .S(rst), 
        .Z(MCInput[56]) );
  MUX2_X1 InputMUX_MUXInst_57_U1 ( .A(Feedback[57]), .B(Input[57]), .S(rst), 
        .Z(MCInput[57]) );
  MUX2_X1 InputMUX_MUXInst_58_U1 ( .A(Feedback[58]), .B(Input[58]), .S(rst), 
        .Z(MCInput[58]) );
  MUX2_X1 InputMUX_MUXInst_59_U1 ( .A(Feedback[59]), .B(Input[59]), .S(rst), 
        .Z(MCInput[59]) );
  MUX2_X1 InputMUX_MUXInst_60_U1 ( .A(Feedback[60]), .B(Input[60]), .S(rst), 
        .Z(MCInput[60]) );
  MUX2_X1 InputMUX_MUXInst_61_U1 ( .A(Feedback[61]), .B(Input[61]), .S(rst), 
        .Z(MCInput[61]) );
  MUX2_X1 InputMUX_MUXInst_62_U1 ( .A(Feedback[62]), .B(Input[62]), .S(rst), 
        .Z(MCInput[62]) );
  MUX2_X1 InputMUX_MUXInst_63_U1 ( .A(Feedback[63]), .B(Input[63]), .S(rst), 
        .Z(MCInput[63]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_0_U3 ( .A(MCInst_XOR_r0_Inst_0_n2), .B(
        MCInst_XOR_r0_Inst_0_n1), .ZN(MCOutput[48]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_0_U2 ( .A(MCOutput[16]), .B(MCOutput[0]), .ZN(
        MCInst_XOR_r0_Inst_0_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_0_U1 ( .A(1'b0), .B(MCInput[48]), .Z(
        MCInst_XOR_r0_Inst_0_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_0_U2 ( .A(MCInst_XOR_r1_Inst_0_n1), .B(
        MCOutput[0]), .ZN(MCOutput[32]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_0_U1 ( .A(1'b0), .B(MCInput[32]), .ZN(
        MCInst_XOR_r1_Inst_0_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U3 ( .A(MCInst_XOR_r0_Inst_1_n2), .B(
        MCInst_XOR_r0_Inst_1_n1), .ZN(MCOutput[49]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U2 ( .A(MCOutput[17]), .B(MCOutput[1]), .ZN(
        MCInst_XOR_r0_Inst_1_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_1_U1 ( .A(1'b0), .B(MCInput[49]), .Z(
        MCInst_XOR_r0_Inst_1_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_1_U2 ( .A(MCInst_XOR_r1_Inst_1_n1), .B(
        MCOutput[1]), .ZN(MCOutput[33]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_1_U1 ( .A(1'b0), .B(MCInput[33]), .ZN(
        MCInst_XOR_r1_Inst_1_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U3 ( .A(MCInst_XOR_r0_Inst_2_n2), .B(
        MCInst_XOR_r0_Inst_2_n1), .ZN(MCOutput[50]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U2 ( .A(MCOutput[18]), .B(MCOutput[2]), .ZN(
        MCInst_XOR_r0_Inst_2_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_2_U1 ( .A(1'b0), .B(MCInput[50]), .Z(
        MCInst_XOR_r0_Inst_2_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_2_U2 ( .A(MCInst_XOR_r1_Inst_2_n1), .B(
        MCOutput[2]), .ZN(MCOutput[34]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_2_U1 ( .A(1'b0), .B(MCInput[34]), .ZN(
        MCInst_XOR_r1_Inst_2_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U3 ( .A(MCInst_XOR_r0_Inst_3_n2), .B(
        MCInst_XOR_r0_Inst_3_n1), .ZN(MCOutput[51]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U2 ( .A(MCOutput[19]), .B(MCOutput[3]), .ZN(
        MCInst_XOR_r0_Inst_3_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_3_U1 ( .A(1'b0), .B(MCInput[51]), .Z(
        MCInst_XOR_r0_Inst_3_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_3_U2 ( .A(MCInst_XOR_r1_Inst_3_n1), .B(
        MCOutput[3]), .ZN(MCOutput[35]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_3_U1 ( .A(1'b0), .B(MCInput[35]), .ZN(
        MCInst_XOR_r1_Inst_3_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U3 ( .A(MCInst_XOR_r0_Inst_4_n2), .B(
        MCInst_XOR_r0_Inst_4_n1), .ZN(MCOutput[52]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U2 ( .A(MCOutput[20]), .B(MCOutput[4]), .ZN(
        MCInst_XOR_r0_Inst_4_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_4_U1 ( .A(1'b0), .B(MCInput[52]), .Z(
        MCInst_XOR_r0_Inst_4_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_4_U2 ( .A(MCInst_XOR_r1_Inst_4_n1), .B(
        MCOutput[4]), .ZN(MCOutput[36]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_4_U1 ( .A(1'b0), .B(MCInput[36]), .ZN(
        MCInst_XOR_r1_Inst_4_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U3 ( .A(MCInst_XOR_r0_Inst_5_n2), .B(
        MCInst_XOR_r0_Inst_5_n1), .ZN(MCOutput[53]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U2 ( .A(MCOutput[21]), .B(MCOutput[5]), .ZN(
        MCInst_XOR_r0_Inst_5_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_5_U1 ( .A(1'b0), .B(MCInput[53]), .Z(
        MCInst_XOR_r0_Inst_5_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_5_U2 ( .A(MCInst_XOR_r1_Inst_5_n1), .B(
        MCOutput[5]), .ZN(MCOutput[37]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_5_U1 ( .A(1'b0), .B(MCInput[37]), .ZN(
        MCInst_XOR_r1_Inst_5_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U3 ( .A(MCInst_XOR_r0_Inst_6_n2), .B(
        MCInst_XOR_r0_Inst_6_n1), .ZN(MCOutput[54]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U2 ( .A(MCOutput[22]), .B(MCOutput[6]), .ZN(
        MCInst_XOR_r0_Inst_6_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_6_U1 ( .A(1'b0), .B(MCInput[54]), .Z(
        MCInst_XOR_r0_Inst_6_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_6_U2 ( .A(MCInst_XOR_r1_Inst_6_n1), .B(
        MCOutput[6]), .ZN(MCOutput[38]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_6_U1 ( .A(1'b0), .B(MCInput[38]), .ZN(
        MCInst_XOR_r1_Inst_6_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U3 ( .A(MCInst_XOR_r0_Inst_7_n2), .B(
        MCInst_XOR_r0_Inst_7_n1), .ZN(MCOutput[55]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U2 ( .A(MCOutput[23]), .B(MCOutput[7]), .ZN(
        MCInst_XOR_r0_Inst_7_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_7_U1 ( .A(1'b0), .B(MCInput[55]), .Z(
        MCInst_XOR_r0_Inst_7_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_7_U2 ( .A(MCInst_XOR_r1_Inst_7_n1), .B(
        MCOutput[7]), .ZN(MCOutput[39]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_7_U1 ( .A(1'b0), .B(MCInput[39]), .ZN(
        MCInst_XOR_r1_Inst_7_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U3 ( .A(MCInst_XOR_r0_Inst_8_n2), .B(
        MCInst_XOR_r0_Inst_8_n1), .ZN(MCOutput[56]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U2 ( .A(MCOutput[24]), .B(MCOutput[8]), .ZN(
        MCInst_XOR_r0_Inst_8_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_8_U1 ( .A(1'b0), .B(MCInput[56]), .Z(
        MCInst_XOR_r0_Inst_8_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_8_U2 ( .A(MCInst_XOR_r1_Inst_8_n1), .B(
        MCOutput[8]), .ZN(MCOutput[40]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_8_U1 ( .A(1'b0), .B(MCInput[40]), .ZN(
        MCInst_XOR_r1_Inst_8_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U3 ( .A(MCInst_XOR_r0_Inst_9_n2), .B(
        MCInst_XOR_r0_Inst_9_n1), .ZN(MCOutput[57]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U2 ( .A(MCOutput[25]), .B(MCOutput[9]), .ZN(
        MCInst_XOR_r0_Inst_9_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_9_U1 ( .A(1'b0), .B(MCInput[57]), .Z(
        MCInst_XOR_r0_Inst_9_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_9_U2 ( .A(MCInst_XOR_r1_Inst_9_n1), .B(
        MCOutput[9]), .ZN(MCOutput[41]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_9_U1 ( .A(1'b0), .B(MCInput[41]), .ZN(
        MCInst_XOR_r1_Inst_9_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U3 ( .A(MCInst_XOR_r0_Inst_10_n2), .B(
        MCInst_XOR_r0_Inst_10_n1), .ZN(MCOutput[58]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U2 ( .A(MCOutput[26]), .B(MCOutput[10]), .ZN(
        MCInst_XOR_r0_Inst_10_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_10_U1 ( .A(1'b0), .B(MCInput[58]), .Z(
        MCInst_XOR_r0_Inst_10_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_10_U2 ( .A(MCInst_XOR_r1_Inst_10_n1), .B(
        MCOutput[10]), .ZN(MCOutput[42]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_10_U1 ( .A(1'b0), .B(MCInput[42]), .ZN(
        MCInst_XOR_r1_Inst_10_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U3 ( .A(MCInst_XOR_r0_Inst_11_n2), .B(
        MCInst_XOR_r0_Inst_11_n1), .ZN(MCOutput[59]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U2 ( .A(MCOutput[27]), .B(MCOutput[11]), .ZN(
        MCInst_XOR_r0_Inst_11_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_11_U1 ( .A(1'b0), .B(MCInput[59]), .Z(
        MCInst_XOR_r0_Inst_11_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_11_U2 ( .A(MCInst_XOR_r1_Inst_11_n1), .B(
        MCOutput[11]), .ZN(MCOutput[43]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_11_U1 ( .A(1'b0), .B(MCInput[43]), .ZN(
        MCInst_XOR_r1_Inst_11_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U3 ( .A(MCInst_XOR_r0_Inst_12_n2), .B(
        MCInst_XOR_r0_Inst_12_n1), .ZN(MCOutput[60]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U2 ( .A(MCOutput[28]), .B(MCOutput[12]), .ZN(
        MCInst_XOR_r0_Inst_12_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_12_U1 ( .A(1'b0), .B(MCInput[60]), .Z(
        MCInst_XOR_r0_Inst_12_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_12_U2 ( .A(MCInst_XOR_r1_Inst_12_n1), .B(
        MCOutput[12]), .ZN(MCOutput[44]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_12_U1 ( .A(1'b0), .B(MCInput[44]), .ZN(
        MCInst_XOR_r1_Inst_12_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U3 ( .A(MCInst_XOR_r0_Inst_13_n2), .B(
        MCInst_XOR_r0_Inst_13_n1), .ZN(MCOutput[61]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U2 ( .A(MCOutput[29]), .B(MCOutput[13]), .ZN(
        MCInst_XOR_r0_Inst_13_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_13_U1 ( .A(1'b0), .B(MCInput[61]), .Z(
        MCInst_XOR_r0_Inst_13_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_13_U2 ( .A(MCInst_XOR_r1_Inst_13_n1), .B(
        MCOutput[13]), .ZN(MCOutput[45]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_13_U1 ( .A(1'b0), .B(MCInput[45]), .ZN(
        MCInst_XOR_r1_Inst_13_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U3 ( .A(MCInst_XOR_r0_Inst_14_n2), .B(
        MCInst_XOR_r0_Inst_14_n1), .ZN(MCOutput[62]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U2 ( .A(MCOutput[30]), .B(MCOutput[14]), .ZN(
        MCInst_XOR_r0_Inst_14_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_14_U1 ( .A(1'b0), .B(MCInput[62]), .Z(
        MCInst_XOR_r0_Inst_14_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_14_U2 ( .A(MCInst_XOR_r1_Inst_14_n1), .B(
        MCOutput[14]), .ZN(MCOutput[46]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_14_U1 ( .A(1'b0), .B(MCInput[46]), .ZN(
        MCInst_XOR_r1_Inst_14_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U3 ( .A(MCInst_XOR_r0_Inst_15_n2), .B(
        MCInst_XOR_r0_Inst_15_n1), .ZN(MCOutput[63]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U2 ( .A(MCOutput[31]), .B(MCOutput[15]), .ZN(
        MCInst_XOR_r0_Inst_15_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_15_U1 ( .A(1'b0), .B(MCInput[63]), .Z(
        MCInst_XOR_r0_Inst_15_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_15_U2 ( .A(MCInst_XOR_r1_Inst_15_n1), .B(
        MCOutput[15]), .ZN(MCOutput[47]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_15_U1 ( .A(1'b0), .B(MCInput[47]), .ZN(
        MCInst_XOR_r1_Inst_15_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_0_U2 ( .A(AddKeyXOR1_XORInst_0_0_n1), .B(
        SelectedKey[48]), .ZN(AddRoundKeyOutput[48]) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_0_U1 ( .A(1'b0), .B(MCOutput[48]), .ZN(
        AddKeyXOR1_XORInst_0_0_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_1_U2 ( .A(AddKeyXOR1_XORInst_0_1_n1), .B(
        SelectedKey[49]), .ZN(AddRoundKeyOutput[49]) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_1_U1 ( .A(1'b0), .B(MCOutput[49]), .ZN(
        AddKeyXOR1_XORInst_0_1_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_2_U2 ( .A(AddKeyXOR1_XORInst_0_2_n1), .B(
        SelectedKey[50]), .ZN(AddRoundKeyOutput[50]) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_2_U1 ( .A(1'b0), .B(MCOutput[50]), .ZN(
        AddKeyXOR1_XORInst_0_2_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_3_U2 ( .A(AddKeyXOR1_XORInst_0_3_n1), .B(
        SelectedKey[51]), .ZN(AddRoundKeyOutput[51]) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_3_U1 ( .A(1'b0), .B(MCOutput[51]), .ZN(
        AddKeyXOR1_XORInst_0_3_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_0_U2 ( .A(AddKeyXOR1_XORInst_1_0_n1), .B(
        SelectedKey[52]), .ZN(AddRoundKeyOutput[52]) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_0_U1 ( .A(1'b0), .B(MCOutput[52]), .ZN(
        AddKeyXOR1_XORInst_1_0_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_1_U2 ( .A(AddKeyXOR1_XORInst_1_1_n1), .B(
        SelectedKey[53]), .ZN(AddRoundKeyOutput[53]) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_1_U1 ( .A(1'b0), .B(MCOutput[53]), .ZN(
        AddKeyXOR1_XORInst_1_1_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_2_U2 ( .A(AddKeyXOR1_XORInst_1_2_n1), .B(
        SelectedKey[54]), .ZN(AddRoundKeyOutput[54]) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_2_U1 ( .A(1'b0), .B(MCOutput[54]), .ZN(
        AddKeyXOR1_XORInst_1_2_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_3_U2 ( .A(AddKeyXOR1_XORInst_1_3_n1), .B(
        SelectedKey[55]), .ZN(AddRoundKeyOutput[55]) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_3_U1 ( .A(1'b0), .B(MCOutput[55]), .ZN(
        AddKeyXOR1_XORInst_1_3_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_0_U2 ( .A(AddKeyXOR1_XORInst_2_0_n1), .B(
        SelectedKey[56]), .ZN(AddRoundKeyOutput[56]) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_0_U1 ( .A(1'b0), .B(MCOutput[56]), .ZN(
        AddKeyXOR1_XORInst_2_0_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_1_U2 ( .A(AddKeyXOR1_XORInst_2_1_n1), .B(
        SelectedKey[57]), .ZN(AddRoundKeyOutput[57]) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_1_U1 ( .A(1'b0), .B(MCOutput[57]), .ZN(
        AddKeyXOR1_XORInst_2_1_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_2_U2 ( .A(AddKeyXOR1_XORInst_2_2_n1), .B(
        SelectedKey[58]), .ZN(AddRoundKeyOutput[58]) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_2_U1 ( .A(1'b0), .B(MCOutput[58]), .ZN(
        AddKeyXOR1_XORInst_2_2_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_3_U2 ( .A(AddKeyXOR1_XORInst_2_3_n1), .B(
        SelectedKey[59]), .ZN(AddRoundKeyOutput[59]) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_3_U1 ( .A(1'b0), .B(MCOutput[59]), .ZN(
        AddKeyXOR1_XORInst_2_3_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_0_U2 ( .A(AddKeyXOR1_XORInst_3_0_n1), .B(
        SelectedKey[60]), .ZN(AddRoundKeyOutput[60]) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_0_U1 ( .A(1'b0), .B(MCOutput[60]), .ZN(
        AddKeyXOR1_XORInst_3_0_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_1_U2 ( .A(AddKeyXOR1_XORInst_3_1_n1), .B(
        SelectedKey[61]), .ZN(AddRoundKeyOutput[61]) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_1_U1 ( .A(1'b0), .B(MCOutput[61]), .ZN(
        AddKeyXOR1_XORInst_3_1_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_2_U2 ( .A(AddKeyXOR1_XORInst_3_2_n1), .B(
        SelectedKey[62]), .ZN(AddRoundKeyOutput[62]) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_2_U1 ( .A(1'b0), .B(MCOutput[62]), .ZN(
        AddKeyXOR1_XORInst_3_2_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_3_U2 ( .A(AddKeyXOR1_XORInst_3_3_n1), .B(
        SelectedKey[63]), .ZN(AddRoundKeyOutput[63]) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_3_U1 ( .A(1'b0), .B(MCOutput[63]), .ZN(
        AddKeyXOR1_XORInst_3_3_n1) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_0_U3 ( .A(AddKeyConstXOR_XORInst_0_0_n2), 
        .B(AddKeyConstXOR_XORInst_0_0_n1), .ZN(AddRoundKeyOutput[40]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_0_U2 ( .A(SelectedKey[40]), .B(
        RoundConstant_0), .ZN(AddKeyConstXOR_XORInst_0_0_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_0_U1 ( .A(1'b0), .B(MCOutput[40]), .Z(
        AddKeyConstXOR_XORInst_0_0_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_1_U3 ( .A(AddKeyConstXOR_XORInst_0_1_n2), 
        .B(AddKeyConstXOR_XORInst_0_1_n1), .ZN(AddRoundKeyOutput[41]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_1_U2 ( .A(SelectedKey[41]), .B(
        FSMUpdate[0]), .ZN(AddKeyConstXOR_XORInst_0_1_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_1_U1 ( .A(1'b0), .B(MCOutput[41]), .Z(
        AddKeyConstXOR_XORInst_0_1_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_2_U3 ( .A(AddKeyConstXOR_XORInst_0_2_n2), 
        .B(AddKeyConstXOR_XORInst_0_2_n1), .ZN(AddRoundKeyOutput[42]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_2_U2 ( .A(SelectedKey[42]), .B(
        FSMUpdate[1]), .ZN(AddKeyConstXOR_XORInst_0_2_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_2_U1 ( .A(1'b0), .B(MCOutput[42]), .Z(
        AddKeyConstXOR_XORInst_0_2_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_3_U3 ( .A(AddKeyConstXOR_XORInst_0_3_n2), 
        .B(AddKeyConstXOR_XORInst_0_3_n1), .ZN(AddRoundKeyOutput[43]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_3_U2 ( .A(SelectedKey[43]), .B(1'b0), .ZN(
        AddKeyConstXOR_XORInst_0_3_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_3_U1 ( .A(1'b0), .B(MCOutput[43]), .Z(
        AddKeyConstXOR_XORInst_0_3_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_0_U3 ( .A(AddKeyConstXOR_XORInst_1_0_n2), 
        .B(AddKeyConstXOR_XORInst_1_0_n1), .ZN(AddRoundKeyOutput[44]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_0_U2 ( .A(SelectedKey[44]), .B(
        RoundConstant_4_), .ZN(AddKeyConstXOR_XORInst_1_0_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_0_U1 ( .A(1'b0), .B(MCOutput[44]), .Z(
        AddKeyConstXOR_XORInst_1_0_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_1_U3 ( .A(AddKeyConstXOR_XORInst_1_1_n2), 
        .B(AddKeyConstXOR_XORInst_1_1_n1), .ZN(AddRoundKeyOutput[45]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_1_U2 ( .A(SelectedKey[45]), .B(
        FSMUpdate[3]), .ZN(AddKeyConstXOR_XORInst_1_1_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_1_U1 ( .A(1'b0), .B(MCOutput[45]), .Z(
        AddKeyConstXOR_XORInst_1_1_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_2_U3 ( .A(AddKeyConstXOR_XORInst_1_2_n2), 
        .B(AddKeyConstXOR_XORInst_1_2_n1), .ZN(AddRoundKeyOutput[46]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_2_U2 ( .A(SelectedKey[46]), .B(
        FSMUpdate[4]), .ZN(AddKeyConstXOR_XORInst_1_2_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_2_U1 ( .A(1'b0), .B(MCOutput[46]), .Z(
        AddKeyConstXOR_XORInst_1_2_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_3_U3 ( .A(AddKeyConstXOR_XORInst_1_3_n2), 
        .B(AddKeyConstXOR_XORInst_1_3_n1), .ZN(AddRoundKeyOutput[47]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_3_U2 ( .A(SelectedKey[47]), .B(
        FSMUpdate[5]), .ZN(AddKeyConstXOR_XORInst_1_3_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_3_U1 ( .A(1'b0), .B(MCOutput[47]), .Z(
        AddKeyConstXOR_XORInst_1_3_n2) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_0_U2 ( .A(AddKeyXOR2_XORInst_0_0_n1), .B(
        SelectedKey[0]), .ZN(AddRoundKeyOutput[0]) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_0_U1 ( .A(1'b0), .B(MCOutput[0]), .ZN(
        AddKeyXOR2_XORInst_0_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_1_U2 ( .A(AddKeyXOR2_XORInst_0_1_n1), .B(
        SelectedKey[1]), .ZN(AddRoundKeyOutput[1]) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_1_U1 ( .A(1'b0), .B(MCOutput[1]), .ZN(
        AddKeyXOR2_XORInst_0_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_2_U2 ( .A(AddKeyXOR2_XORInst_0_2_n1), .B(
        SelectedKey[2]), .ZN(AddRoundKeyOutput[2]) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_2_U1 ( .A(1'b0), .B(MCOutput[2]), .ZN(
        AddKeyXOR2_XORInst_0_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_3_U2 ( .A(AddKeyXOR2_XORInst_0_3_n1), .B(
        SelectedKey[3]), .ZN(AddRoundKeyOutput[3]) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_3_U1 ( .A(1'b0), .B(MCOutput[3]), .ZN(
        AddKeyXOR2_XORInst_0_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_0_U2 ( .A(AddKeyXOR2_XORInst_1_0_n1), .B(
        SelectedKey[4]), .ZN(AddRoundKeyOutput[4]) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_0_U1 ( .A(1'b0), .B(MCOutput[4]), .ZN(
        AddKeyXOR2_XORInst_1_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_1_U2 ( .A(AddKeyXOR2_XORInst_1_1_n1), .B(
        SelectedKey[5]), .ZN(AddRoundKeyOutput[5]) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_1_U1 ( .A(1'b0), .B(MCOutput[5]), .ZN(
        AddKeyXOR2_XORInst_1_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_2_U2 ( .A(AddKeyXOR2_XORInst_1_2_n1), .B(
        SelectedKey[6]), .ZN(AddRoundKeyOutput[6]) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_2_U1 ( .A(1'b0), .B(MCOutput[6]), .ZN(
        AddKeyXOR2_XORInst_1_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_3_U2 ( .A(AddKeyXOR2_XORInst_1_3_n1), .B(
        SelectedKey[7]), .ZN(AddRoundKeyOutput[7]) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_3_U1 ( .A(1'b0), .B(MCOutput[7]), .ZN(
        AddKeyXOR2_XORInst_1_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_0_U2 ( .A(AddKeyXOR2_XORInst_2_0_n1), .B(
        SelectedKey[8]), .ZN(AddRoundKeyOutput[8]) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_0_U1 ( .A(1'b0), .B(MCOutput[8]), .ZN(
        AddKeyXOR2_XORInst_2_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_1_U2 ( .A(AddKeyXOR2_XORInst_2_1_n1), .B(
        SelectedKey[9]), .ZN(AddRoundKeyOutput[9]) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_1_U1 ( .A(1'b0), .B(MCOutput[9]), .ZN(
        AddKeyXOR2_XORInst_2_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_2_U2 ( .A(AddKeyXOR2_XORInst_2_2_n1), .B(
        SelectedKey[10]), .ZN(AddRoundKeyOutput[10]) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_2_U1 ( .A(1'b0), .B(MCOutput[10]), .ZN(
        AddKeyXOR2_XORInst_2_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_3_U2 ( .A(AddKeyXOR2_XORInst_2_3_n1), .B(
        SelectedKey[11]), .ZN(AddRoundKeyOutput[11]) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_3_U1 ( .A(1'b0), .B(MCOutput[11]), .ZN(
        AddKeyXOR2_XORInst_2_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_0_U2 ( .A(AddKeyXOR2_XORInst_3_0_n1), .B(
        SelectedKey[12]), .ZN(AddRoundKeyOutput[12]) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_0_U1 ( .A(1'b0), .B(MCOutput[12]), .ZN(
        AddKeyXOR2_XORInst_3_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_1_U2 ( .A(AddKeyXOR2_XORInst_3_1_n1), .B(
        SelectedKey[13]), .ZN(AddRoundKeyOutput[13]) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_1_U1 ( .A(1'b0), .B(MCOutput[13]), .ZN(
        AddKeyXOR2_XORInst_3_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_2_U2 ( .A(AddKeyXOR2_XORInst_3_2_n1), .B(
        SelectedKey[14]), .ZN(AddRoundKeyOutput[14]) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_2_U1 ( .A(1'b0), .B(MCOutput[14]), .ZN(
        AddKeyXOR2_XORInst_3_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_3_U2 ( .A(AddKeyXOR2_XORInst_3_3_n1), .B(
        SelectedKey[15]), .ZN(AddRoundKeyOutput[15]) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_3_U1 ( .A(1'b0), .B(MCOutput[15]), .ZN(
        AddKeyXOR2_XORInst_3_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_0_U2 ( .A(AddKeyXOR2_XORInst_4_0_n1), .B(
        SelectedKey[16]), .ZN(AddRoundKeyOutput[16]) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_0_U1 ( .A(1'b0), .B(MCOutput[16]), .ZN(
        AddKeyXOR2_XORInst_4_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_1_U2 ( .A(AddKeyXOR2_XORInst_4_1_n1), .B(
        SelectedKey[17]), .ZN(AddRoundKeyOutput[17]) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_1_U1 ( .A(1'b0), .B(MCOutput[17]), .ZN(
        AddKeyXOR2_XORInst_4_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_2_U2 ( .A(AddKeyXOR2_XORInst_4_2_n1), .B(
        SelectedKey[18]), .ZN(AddRoundKeyOutput[18]) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_2_U1 ( .A(1'b0), .B(MCOutput[18]), .ZN(
        AddKeyXOR2_XORInst_4_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_3_U2 ( .A(AddKeyXOR2_XORInst_4_3_n1), .B(
        SelectedKey[19]), .ZN(AddRoundKeyOutput[19]) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_3_U1 ( .A(1'b0), .B(MCOutput[19]), .ZN(
        AddKeyXOR2_XORInst_4_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_0_U2 ( .A(AddKeyXOR2_XORInst_5_0_n1), .B(
        SelectedKey[20]), .ZN(AddRoundKeyOutput[20]) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_0_U1 ( .A(1'b0), .B(MCOutput[20]), .ZN(
        AddKeyXOR2_XORInst_5_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_1_U2 ( .A(AddKeyXOR2_XORInst_5_1_n1), .B(
        SelectedKey[21]), .ZN(AddRoundKeyOutput[21]) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_1_U1 ( .A(1'b0), .B(MCOutput[21]), .ZN(
        AddKeyXOR2_XORInst_5_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_2_U2 ( .A(AddKeyXOR2_XORInst_5_2_n1), .B(
        SelectedKey[22]), .ZN(AddRoundKeyOutput[22]) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_2_U1 ( .A(1'b0), .B(MCOutput[22]), .ZN(
        AddKeyXOR2_XORInst_5_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_3_U2 ( .A(AddKeyXOR2_XORInst_5_3_n1), .B(
        SelectedKey[23]), .ZN(AddRoundKeyOutput[23]) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_3_U1 ( .A(1'b0), .B(MCOutput[23]), .ZN(
        AddKeyXOR2_XORInst_5_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_0_U2 ( .A(AddKeyXOR2_XORInst_6_0_n1), .B(
        SelectedKey[24]), .ZN(AddRoundKeyOutput[24]) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_0_U1 ( .A(1'b0), .B(MCOutput[24]), .ZN(
        AddKeyXOR2_XORInst_6_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_1_U2 ( .A(AddKeyXOR2_XORInst_6_1_n1), .B(
        SelectedKey[25]), .ZN(AddRoundKeyOutput[25]) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_1_U1 ( .A(1'b0), .B(MCOutput[25]), .ZN(
        AddKeyXOR2_XORInst_6_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_2_U2 ( .A(AddKeyXOR2_XORInst_6_2_n1), .B(
        SelectedKey[26]), .ZN(AddRoundKeyOutput[26]) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_2_U1 ( .A(1'b0), .B(MCOutput[26]), .ZN(
        AddKeyXOR2_XORInst_6_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_3_U2 ( .A(AddKeyXOR2_XORInst_6_3_n1), .B(
        SelectedKey[27]), .ZN(AddRoundKeyOutput[27]) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_3_U1 ( .A(1'b0), .B(MCOutput[27]), .ZN(
        AddKeyXOR2_XORInst_6_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_0_U2 ( .A(AddKeyXOR2_XORInst_7_0_n1), .B(
        SelectedKey[28]), .ZN(AddRoundKeyOutput[28]) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_0_U1 ( .A(1'b0), .B(MCOutput[28]), .ZN(
        AddKeyXOR2_XORInst_7_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_1_U2 ( .A(AddKeyXOR2_XORInst_7_1_n1), .B(
        SelectedKey[29]), .ZN(AddRoundKeyOutput[29]) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_1_U1 ( .A(1'b0), .B(MCOutput[29]), .ZN(
        AddKeyXOR2_XORInst_7_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_2_U2 ( .A(AddKeyXOR2_XORInst_7_2_n1), .B(
        SelectedKey[30]), .ZN(AddRoundKeyOutput[30]) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_2_U1 ( .A(1'b0), .B(MCOutput[30]), .ZN(
        AddKeyXOR2_XORInst_7_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_3_U2 ( .A(AddKeyXOR2_XORInst_7_3_n1), .B(
        SelectedKey[31]), .ZN(AddRoundKeyOutput[31]) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_3_U1 ( .A(1'b0), .B(MCOutput[31]), .ZN(
        AddKeyXOR2_XORInst_7_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_0_U2 ( .A(AddKeyXOR2_XORInst_8_0_n1), .B(
        SelectedKey[32]), .ZN(AddRoundKeyOutput[32]) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_0_U1 ( .A(1'b0), .B(MCOutput[32]), .ZN(
        AddKeyXOR2_XORInst_8_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_1_U2 ( .A(AddKeyXOR2_XORInst_8_1_n1), .B(
        SelectedKey[33]), .ZN(AddRoundKeyOutput[33]) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_1_U1 ( .A(1'b0), .B(MCOutput[33]), .ZN(
        AddKeyXOR2_XORInst_8_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_2_U2 ( .A(AddKeyXOR2_XORInst_8_2_n1), .B(
        SelectedKey[34]), .ZN(AddRoundKeyOutput[34]) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_2_U1 ( .A(1'b0), .B(MCOutput[34]), .ZN(
        AddKeyXOR2_XORInst_8_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_3_U2 ( .A(AddKeyXOR2_XORInst_8_3_n1), .B(
        SelectedKey[35]), .ZN(AddRoundKeyOutput[35]) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_3_U1 ( .A(1'b0), .B(MCOutput[35]), .ZN(
        AddKeyXOR2_XORInst_8_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_0_U2 ( .A(AddKeyXOR2_XORInst_9_0_n1), .B(
        SelectedKey[36]), .ZN(AddRoundKeyOutput[36]) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_0_U1 ( .A(1'b0), .B(MCOutput[36]), .ZN(
        AddKeyXOR2_XORInst_9_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_1_U2 ( .A(AddKeyXOR2_XORInst_9_1_n1), .B(
        SelectedKey[37]), .ZN(AddRoundKeyOutput[37]) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_1_U1 ( .A(1'b0), .B(MCOutput[37]), .ZN(
        AddKeyXOR2_XORInst_9_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_2_U2 ( .A(AddKeyXOR2_XORInst_9_2_n1), .B(
        SelectedKey[38]), .ZN(AddRoundKeyOutput[38]) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_2_U1 ( .A(1'b0), .B(MCOutput[38]), .ZN(
        AddKeyXOR2_XORInst_9_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_3_U2 ( .A(AddKeyXOR2_XORInst_9_3_n1), .B(
        SelectedKey[39]), .ZN(AddRoundKeyOutput[39]) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_3_U1 ( .A(1'b0), .B(MCOutput[39]), .ZN(
        AddKeyXOR2_XORInst_9_3_n1) );
  DFF_X1 StateReg_s_current_state_reg_0_ ( .D(AddRoundKeyOutput[0]), .CK(clk), 
        .Q(PermutationOutput[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1_ ( .D(AddRoundKeyOutput[1]), .CK(clk), 
        .Q(PermutationOutput[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2_ ( .D(AddRoundKeyOutput[2]), .CK(clk), 
        .Q(PermutationOutput[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3_ ( .D(AddRoundKeyOutput[3]), .CK(clk), 
        .Q(PermutationOutput[63]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4_ ( .D(AddRoundKeyOutput[4]), .CK(clk), 
        .Q(PermutationOutput[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5_ ( .D(AddRoundKeyOutput[5]), .CK(clk), 
        .Q(PermutationOutput[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6_ ( .D(AddRoundKeyOutput[6]), .CK(clk), 
        .Q(PermutationOutput[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7_ ( .D(AddRoundKeyOutput[7]), .CK(clk), 
        .Q(PermutationOutput[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8_ ( .D(AddRoundKeyOutput[8]), .CK(clk), 
        .Q(PermutationOutput[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9_ ( .D(AddRoundKeyOutput[9]), .CK(clk), 
        .Q(PermutationOutput[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10_ ( .D(AddRoundKeyOutput[10]), .CK(clk), .Q(PermutationOutput[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11_ ( .D(AddRoundKeyOutput[11]), .CK(clk), .Q(PermutationOutput[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12_ ( .D(AddRoundKeyOutput[12]), .CK(clk), .Q(PermutationOutput[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13_ ( .D(AddRoundKeyOutput[13]), .CK(clk), .Q(PermutationOutput[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14_ ( .D(AddRoundKeyOutput[14]), .CK(clk), .Q(PermutationOutput[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15_ ( .D(AddRoundKeyOutput[15]), .CK(clk), .Q(PermutationOutput[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16_ ( .D(AddRoundKeyOutput[16]), .CK(clk), .Q(PermutationOutput[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17_ ( .D(AddRoundKeyOutput[17]), .CK(clk), .Q(PermutationOutput[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18_ ( .D(AddRoundKeyOutput[18]), .CK(clk), .Q(PermutationOutput[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19_ ( .D(AddRoundKeyOutput[19]), .CK(clk), .Q(PermutationOutput[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20_ ( .D(AddRoundKeyOutput[20]), .CK(clk), .Q(PermutationOutput[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21_ ( .D(AddRoundKeyOutput[21]), .CK(clk), .Q(PermutationOutput[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22_ ( .D(AddRoundKeyOutput[22]), .CK(clk), .Q(PermutationOutput[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23_ ( .D(AddRoundKeyOutput[23]), .CK(clk), .Q(PermutationOutput[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24_ ( .D(AddRoundKeyOutput[24]), .CK(clk), .Q(PermutationOutput[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25_ ( .D(AddRoundKeyOutput[25]), .CK(clk), .Q(PermutationOutput[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26_ ( .D(AddRoundKeyOutput[26]), .CK(clk), .Q(PermutationOutput[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27_ ( .D(AddRoundKeyOutput[27]), .CK(clk), .Q(PermutationOutput[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28_ ( .D(AddRoundKeyOutput[28]), .CK(clk), .Q(PermutationOutput[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29_ ( .D(AddRoundKeyOutput[29]), .CK(clk), .Q(PermutationOutput[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30_ ( .D(AddRoundKeyOutput[30]), .CK(clk), .Q(PermutationOutput[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31_ ( .D(AddRoundKeyOutput[31]), .CK(clk), .Q(PermutationOutput[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32_ ( .D(AddRoundKeyOutput[32]), .CK(clk), .Q(PermutationOutput[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33_ ( .D(AddRoundKeyOutput[33]), .CK(clk), .Q(PermutationOutput[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34_ ( .D(AddRoundKeyOutput[34]), .CK(clk), .Q(PermutationOutput[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35_ ( .D(AddRoundKeyOutput[35]), .CK(clk), .Q(PermutationOutput[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36_ ( .D(AddRoundKeyOutput[36]), .CK(clk), .Q(PermutationOutput[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37_ ( .D(AddRoundKeyOutput[37]), .CK(clk), .Q(PermutationOutput[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38_ ( .D(AddRoundKeyOutput[38]), .CK(clk), .Q(PermutationOutput[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39_ ( .D(AddRoundKeyOutput[39]), .CK(clk), .Q(PermutationOutput[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40_ ( .D(AddRoundKeyOutput[40]), .CK(clk), .Q(PermutationOutput[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41_ ( .D(AddRoundKeyOutput[41]), .CK(clk), .Q(PermutationOutput[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42_ ( .D(AddRoundKeyOutput[42]), .CK(clk), .Q(PermutationOutput[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43_ ( .D(AddRoundKeyOutput[43]), .CK(clk), .Q(PermutationOutput[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44_ ( .D(AddRoundKeyOutput[44]), .CK(clk), .Q(PermutationOutput[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45_ ( .D(AddRoundKeyOutput[45]), .CK(clk), .Q(PermutationOutput[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46_ ( .D(AddRoundKeyOutput[46]), .CK(clk), .Q(PermutationOutput[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47_ ( .D(AddRoundKeyOutput[47]), .CK(clk), .Q(PermutationOutput[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48_ ( .D(AddRoundKeyOutput[48]), .CK(clk), .Q(PermutationOutput[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49_ ( .D(AddRoundKeyOutput[49]), .CK(clk), .Q(PermutationOutput[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50_ ( .D(AddRoundKeyOutput[50]), .CK(clk), .Q(PermutationOutput[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51_ ( .D(AddRoundKeyOutput[51]), .CK(clk), .Q(PermutationOutput[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52_ ( .D(AddRoundKeyOutput[52]), .CK(clk), .Q(PermutationOutput[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53_ ( .D(AddRoundKeyOutput[53]), .CK(clk), .Q(PermutationOutput[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54_ ( .D(AddRoundKeyOutput[54]), .CK(clk), .Q(PermutationOutput[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55_ ( .D(AddRoundKeyOutput[55]), .CK(clk), .Q(PermutationOutput[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56_ ( .D(AddRoundKeyOutput[56]), .CK(clk), .Q(PermutationOutput[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57_ ( .D(AddRoundKeyOutput[57]), .CK(clk), .Q(PermutationOutput[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58_ ( .D(AddRoundKeyOutput[58]), .CK(clk), .Q(PermutationOutput[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59_ ( .D(AddRoundKeyOutput[59]), .CK(clk), .Q(PermutationOutput[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60_ ( .D(AddRoundKeyOutput[60]), .CK(clk), .Q(PermutationOutput[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61_ ( .D(AddRoundKeyOutput[61]), .CK(clk), .Q(PermutationOutput[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62_ ( .D(AddRoundKeyOutput[62]), .CK(clk), .Q(PermutationOutput[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63_ ( .D(AddRoundKeyOutput[63]), .CK(clk), .Q(PermutationOutput[3]), .QN() );
  AOI21_X1 SubCellInst_LFInst_0_LFInst_0_U2 ( .B1(PermutationOutput[3]), .B2(
        PermutationOutput[2]), .A(SubCellInst_LFInst_0_LFInst_0_n1), .ZN(
        Feedback[0]) );
  AOI221_X1 SubCellInst_LFInst_0_LFInst_0_U1 ( .B1(PermutationOutput[2]), .B2(
        PermutationOutput[0]), .C1(PermutationOutput[3]), .C2(
        PermutationOutput[0]), .A(PermutationOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_0_LFInst_1_U3 ( .B1(PermutationOutput[3]), .B2(
        SubCellInst_LFInst_0_LFInst_1_n2), .A(SubCellInst_LFInst_0_LFInst_1_n1), .ZN(Feedback[1]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U2 ( .A1(PermutationOutput[0]), .A2(
        PermutationOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_1_U1 ( .A1(PermutationOutput[0]), .A2(
        PermutationOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_0_LFInst_2_U2 ( .B1(PermutationOutput[3]), .B2(
        PermutationOutput[0]), .A(SubCellInst_LFInst_0_LFInst_2_n1), .ZN(
        Feedback[2]) );
  OAI221_X1 SubCellInst_LFInst_0_LFInst_2_U1 ( .B1(PermutationOutput[2]), .B2(
        PermutationOutput[3]), .C1(PermutationOutput[2]), .C2(
        PermutationOutput[0]), .A(PermutationOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_0_LFInst_3_U1 ( .A1(PermutationOutput[1]), .A2(
        PermutationOutput[3]), .B1(PermutationOutput[1]), .B2(
        PermutationOutput[0]), .C1(PermutationOutput[3]), .C2(
        PermutationOutput[2]), .ZN(Feedback[3]) );
  AOI21_X1 SubCellInst_LFInst_1_LFInst_0_U2 ( .B1(PermutationOutput[7]), .B2(
        PermutationOutput[6]), .A(SubCellInst_LFInst_1_LFInst_0_n1), .ZN(
        Feedback[4]) );
  AOI221_X1 SubCellInst_LFInst_1_LFInst_0_U1 ( .B1(PermutationOutput[6]), .B2(
        PermutationOutput[4]), .C1(PermutationOutput[7]), .C2(
        PermutationOutput[4]), .A(PermutationOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_1_LFInst_1_U3 ( .B1(PermutationOutput[7]), .B2(
        SubCellInst_LFInst_1_LFInst_1_n2), .A(SubCellInst_LFInst_1_LFInst_1_n1), .ZN(Feedback[5]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U2 ( .A1(PermutationOutput[4]), .A2(
        PermutationOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_1_U1 ( .A1(PermutationOutput[4]), .A2(
        PermutationOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_1_LFInst_2_U2 ( .B1(PermutationOutput[7]), .B2(
        PermutationOutput[4]), .A(SubCellInst_LFInst_1_LFInst_2_n1), .ZN(
        Feedback[6]) );
  OAI221_X1 SubCellInst_LFInst_1_LFInst_2_U1 ( .B1(PermutationOutput[6]), .B2(
        PermutationOutput[7]), .C1(PermutationOutput[6]), .C2(
        PermutationOutput[4]), .A(PermutationOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_1_LFInst_3_U1 ( .A1(PermutationOutput[5]), .A2(
        PermutationOutput[7]), .B1(PermutationOutput[5]), .B2(
        PermutationOutput[4]), .C1(PermutationOutput[7]), .C2(
        PermutationOutput[6]), .ZN(Feedback[7]) );
  AOI21_X1 SubCellInst_LFInst_2_LFInst_0_U2 ( .B1(PermutationOutput[11]), .B2(
        PermutationOutput[10]), .A(SubCellInst_LFInst_2_LFInst_0_n1), .ZN(
        Feedback[8]) );
  AOI221_X1 SubCellInst_LFInst_2_LFInst_0_U1 ( .B1(PermutationOutput[10]), 
        .B2(PermutationOutput[8]), .C1(PermutationOutput[11]), .C2(
        PermutationOutput[8]), .A(PermutationOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_2_LFInst_1_U3 ( .B1(PermutationOutput[11]), .B2(
        SubCellInst_LFInst_2_LFInst_1_n2), .A(SubCellInst_LFInst_2_LFInst_1_n1), .ZN(Feedback[9]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U2 ( .A1(PermutationOutput[8]), .A2(
        PermutationOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_1_U1 ( .A1(PermutationOutput[8]), .A2(
        PermutationOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_2_LFInst_2_U2 ( .B1(PermutationOutput[11]), .B2(
        PermutationOutput[8]), .A(SubCellInst_LFInst_2_LFInst_2_n1), .ZN(
        Feedback[10]) );
  OAI221_X1 SubCellInst_LFInst_2_LFInst_2_U1 ( .B1(PermutationOutput[10]), 
        .B2(PermutationOutput[11]), .C1(PermutationOutput[10]), .C2(
        PermutationOutput[8]), .A(PermutationOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_2_LFInst_3_U1 ( .A1(PermutationOutput[9]), .A2(
        PermutationOutput[11]), .B1(PermutationOutput[9]), .B2(
        PermutationOutput[8]), .C1(PermutationOutput[11]), .C2(
        PermutationOutput[10]), .ZN(Feedback[11]) );
  AOI21_X1 SubCellInst_LFInst_3_LFInst_0_U2 ( .B1(PermutationOutput[15]), .B2(
        PermutationOutput[14]), .A(SubCellInst_LFInst_3_LFInst_0_n1), .ZN(
        Feedback[12]) );
  AOI221_X1 SubCellInst_LFInst_3_LFInst_0_U1 ( .B1(PermutationOutput[14]), 
        .B2(PermutationOutput[12]), .C1(PermutationOutput[15]), .C2(
        PermutationOutput[12]), .A(PermutationOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_3_LFInst_1_U3 ( .B1(PermutationOutput[15]), .B2(
        SubCellInst_LFInst_3_LFInst_1_n2), .A(SubCellInst_LFInst_3_LFInst_1_n1), .ZN(Feedback[13]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U2 ( .A1(PermutationOutput[12]), .A2(
        PermutationOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_1_U1 ( .A1(PermutationOutput[12]), .A2(
        PermutationOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_3_LFInst_2_U2 ( .B1(PermutationOutput[15]), .B2(
        PermutationOutput[12]), .A(SubCellInst_LFInst_3_LFInst_2_n1), .ZN(
        Feedback[14]) );
  OAI221_X1 SubCellInst_LFInst_3_LFInst_2_U1 ( .B1(PermutationOutput[14]), 
        .B2(PermutationOutput[15]), .C1(PermutationOutput[14]), .C2(
        PermutationOutput[12]), .A(PermutationOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_3_LFInst_3_U1 ( .A1(PermutationOutput[13]), 
        .A2(PermutationOutput[15]), .B1(PermutationOutput[13]), .B2(
        PermutationOutput[12]), .C1(PermutationOutput[15]), .C2(
        PermutationOutput[14]), .ZN(Feedback[15]) );
  AOI21_X1 SubCellInst_LFInst_4_LFInst_0_U2 ( .B1(PermutationOutput[19]), .B2(
        PermutationOutput[18]), .A(SubCellInst_LFInst_4_LFInst_0_n1), .ZN(
        Feedback[16]) );
  AOI221_X1 SubCellInst_LFInst_4_LFInst_0_U1 ( .B1(PermutationOutput[18]), 
        .B2(PermutationOutput[16]), .C1(PermutationOutput[19]), .C2(
        PermutationOutput[16]), .A(PermutationOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_4_LFInst_1_U3 ( .B1(PermutationOutput[19]), .B2(
        SubCellInst_LFInst_4_LFInst_1_n2), .A(SubCellInst_LFInst_4_LFInst_1_n1), .ZN(Feedback[17]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U2 ( .A1(PermutationOutput[16]), .A2(
        PermutationOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_1_U1 ( .A1(PermutationOutput[16]), .A2(
        PermutationOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_4_LFInst_2_U2 ( .B1(PermutationOutput[19]), .B2(
        PermutationOutput[16]), .A(SubCellInst_LFInst_4_LFInst_2_n1), .ZN(
        Feedback[18]) );
  OAI221_X1 SubCellInst_LFInst_4_LFInst_2_U1 ( .B1(PermutationOutput[18]), 
        .B2(PermutationOutput[19]), .C1(PermutationOutput[18]), .C2(
        PermutationOutput[16]), .A(PermutationOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_4_LFInst_3_U1 ( .A1(PermutationOutput[17]), 
        .A2(PermutationOutput[19]), .B1(PermutationOutput[17]), .B2(
        PermutationOutput[16]), .C1(PermutationOutput[19]), .C2(
        PermutationOutput[18]), .ZN(Feedback[19]) );
  AOI21_X1 SubCellInst_LFInst_5_LFInst_0_U2 ( .B1(PermutationOutput[23]), .B2(
        PermutationOutput[22]), .A(SubCellInst_LFInst_5_LFInst_0_n1), .ZN(
        Feedback[20]) );
  AOI221_X1 SubCellInst_LFInst_5_LFInst_0_U1 ( .B1(PermutationOutput[22]), 
        .B2(PermutationOutput[20]), .C1(PermutationOutput[23]), .C2(
        PermutationOutput[20]), .A(PermutationOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_5_LFInst_1_U3 ( .B1(PermutationOutput[23]), .B2(
        SubCellInst_LFInst_5_LFInst_1_n2), .A(SubCellInst_LFInst_5_LFInst_1_n1), .ZN(Feedback[21]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U2 ( .A1(PermutationOutput[20]), .A2(
        PermutationOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_1_U1 ( .A1(PermutationOutput[20]), .A2(
        PermutationOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_5_LFInst_2_U2 ( .B1(PermutationOutput[23]), .B2(
        PermutationOutput[20]), .A(SubCellInst_LFInst_5_LFInst_2_n1), .ZN(
        Feedback[22]) );
  OAI221_X1 SubCellInst_LFInst_5_LFInst_2_U1 ( .B1(PermutationOutput[22]), 
        .B2(PermutationOutput[23]), .C1(PermutationOutput[22]), .C2(
        PermutationOutput[20]), .A(PermutationOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_5_LFInst_3_U1 ( .A1(PermutationOutput[21]), 
        .A2(PermutationOutput[23]), .B1(PermutationOutput[21]), .B2(
        PermutationOutput[20]), .C1(PermutationOutput[23]), .C2(
        PermutationOutput[22]), .ZN(Feedback[23]) );
  AOI21_X1 SubCellInst_LFInst_6_LFInst_0_U2 ( .B1(PermutationOutput[27]), .B2(
        PermutationOutput[26]), .A(SubCellInst_LFInst_6_LFInst_0_n1), .ZN(
        Feedback[24]) );
  AOI221_X1 SubCellInst_LFInst_6_LFInst_0_U1 ( .B1(PermutationOutput[26]), 
        .B2(PermutationOutput[24]), .C1(PermutationOutput[27]), .C2(
        PermutationOutput[24]), .A(PermutationOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_6_LFInst_1_U3 ( .B1(PermutationOutput[27]), .B2(
        SubCellInst_LFInst_6_LFInst_1_n2), .A(SubCellInst_LFInst_6_LFInst_1_n1), .ZN(Feedback[25]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U2 ( .A1(PermutationOutput[24]), .A2(
        PermutationOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_1_U1 ( .A1(PermutationOutput[24]), .A2(
        PermutationOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_6_LFInst_2_U2 ( .B1(PermutationOutput[27]), .B2(
        PermutationOutput[24]), .A(SubCellInst_LFInst_6_LFInst_2_n1), .ZN(
        Feedback[26]) );
  OAI221_X1 SubCellInst_LFInst_6_LFInst_2_U1 ( .B1(PermutationOutput[26]), 
        .B2(PermutationOutput[27]), .C1(PermutationOutput[26]), .C2(
        PermutationOutput[24]), .A(PermutationOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_6_LFInst_3_U1 ( .A1(PermutationOutput[25]), 
        .A2(PermutationOutput[27]), .B1(PermutationOutput[25]), .B2(
        PermutationOutput[24]), .C1(PermutationOutput[27]), .C2(
        PermutationOutput[26]), .ZN(Feedback[27]) );
  AOI21_X1 SubCellInst_LFInst_7_LFInst_0_U2 ( .B1(PermutationOutput[31]), .B2(
        PermutationOutput[30]), .A(SubCellInst_LFInst_7_LFInst_0_n1), .ZN(
        Feedback[28]) );
  AOI221_X1 SubCellInst_LFInst_7_LFInst_0_U1 ( .B1(PermutationOutput[30]), 
        .B2(PermutationOutput[28]), .C1(PermutationOutput[31]), .C2(
        PermutationOutput[28]), .A(PermutationOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_7_LFInst_1_U3 ( .B1(PermutationOutput[31]), .B2(
        SubCellInst_LFInst_7_LFInst_1_n2), .A(SubCellInst_LFInst_7_LFInst_1_n1), .ZN(Feedback[29]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U2 ( .A1(PermutationOutput[28]), .A2(
        PermutationOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_1_U1 ( .A1(PermutationOutput[28]), .A2(
        PermutationOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_7_LFInst_2_U2 ( .B1(PermutationOutput[31]), .B2(
        PermutationOutput[28]), .A(SubCellInst_LFInst_7_LFInst_2_n1), .ZN(
        Feedback[30]) );
  OAI221_X1 SubCellInst_LFInst_7_LFInst_2_U1 ( .B1(PermutationOutput[30]), 
        .B2(PermutationOutput[31]), .C1(PermutationOutput[30]), .C2(
        PermutationOutput[28]), .A(PermutationOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_7_LFInst_3_U1 ( .A1(PermutationOutput[29]), 
        .A2(PermutationOutput[31]), .B1(PermutationOutput[29]), .B2(
        PermutationOutput[28]), .C1(PermutationOutput[31]), .C2(
        PermutationOutput[30]), .ZN(Feedback[31]) );
  AOI21_X1 SubCellInst_LFInst_8_LFInst_0_U2 ( .B1(PermutationOutput[35]), .B2(
        PermutationOutput[34]), .A(SubCellInst_LFInst_8_LFInst_0_n1), .ZN(
        Feedback[32]) );
  AOI221_X1 SubCellInst_LFInst_8_LFInst_0_U1 ( .B1(PermutationOutput[34]), 
        .B2(PermutationOutput[32]), .C1(PermutationOutput[35]), .C2(
        PermutationOutput[32]), .A(PermutationOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_8_LFInst_1_U3 ( .B1(PermutationOutput[35]), .B2(
        SubCellInst_LFInst_8_LFInst_1_n2), .A(SubCellInst_LFInst_8_LFInst_1_n1), .ZN(Feedback[33]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U2 ( .A1(PermutationOutput[32]), .A2(
        PermutationOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_1_U1 ( .A1(PermutationOutput[32]), .A2(
        PermutationOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_8_LFInst_2_U2 ( .B1(PermutationOutput[35]), .B2(
        PermutationOutput[32]), .A(SubCellInst_LFInst_8_LFInst_2_n1), .ZN(
        Feedback[34]) );
  OAI221_X1 SubCellInst_LFInst_8_LFInst_2_U1 ( .B1(PermutationOutput[34]), 
        .B2(PermutationOutput[35]), .C1(PermutationOutput[34]), .C2(
        PermutationOutput[32]), .A(PermutationOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_8_LFInst_3_U1 ( .A1(PermutationOutput[33]), 
        .A2(PermutationOutput[35]), .B1(PermutationOutput[33]), .B2(
        PermutationOutput[32]), .C1(PermutationOutput[35]), .C2(
        PermutationOutput[34]), .ZN(Feedback[35]) );
  AOI21_X1 SubCellInst_LFInst_9_LFInst_0_U2 ( .B1(PermutationOutput[39]), .B2(
        PermutationOutput[38]), .A(SubCellInst_LFInst_9_LFInst_0_n1), .ZN(
        Feedback[36]) );
  AOI221_X1 SubCellInst_LFInst_9_LFInst_0_U1 ( .B1(PermutationOutput[38]), 
        .B2(PermutationOutput[36]), .C1(PermutationOutput[39]), .C2(
        PermutationOutput[36]), .A(PermutationOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_9_LFInst_1_U3 ( .B1(PermutationOutput[39]), .B2(
        SubCellInst_LFInst_9_LFInst_1_n2), .A(SubCellInst_LFInst_9_LFInst_1_n1), .ZN(Feedback[37]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U2 ( .A1(PermutationOutput[36]), .A2(
        PermutationOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_1_U1 ( .A1(PermutationOutput[36]), .A2(
        PermutationOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_9_LFInst_2_U2 ( .B1(PermutationOutput[39]), .B2(
        PermutationOutput[36]), .A(SubCellInst_LFInst_9_LFInst_2_n1), .ZN(
        Feedback[38]) );
  OAI221_X1 SubCellInst_LFInst_9_LFInst_2_U1 ( .B1(PermutationOutput[38]), 
        .B2(PermutationOutput[39]), .C1(PermutationOutput[38]), .C2(
        PermutationOutput[36]), .A(PermutationOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_9_LFInst_3_U1 ( .A1(PermutationOutput[37]), 
        .A2(PermutationOutput[39]), .B1(PermutationOutput[37]), .B2(
        PermutationOutput[36]), .C1(PermutationOutput[39]), .C2(
        PermutationOutput[38]), .ZN(Feedback[39]) );
  AOI21_X1 SubCellInst_LFInst_10_LFInst_0_U2 ( .B1(PermutationOutput[43]), 
        .B2(PermutationOutput[42]), .A(SubCellInst_LFInst_10_LFInst_0_n1), 
        .ZN(Feedback[40]) );
  AOI221_X1 SubCellInst_LFInst_10_LFInst_0_U1 ( .B1(PermutationOutput[42]), 
        .B2(PermutationOutput[40]), .C1(PermutationOutput[43]), .C2(
        PermutationOutput[40]), .A(PermutationOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_10_LFInst_1_U3 ( .B1(PermutationOutput[43]), 
        .B2(SubCellInst_LFInst_10_LFInst_1_n2), .A(
        SubCellInst_LFInst_10_LFInst_1_n1), .ZN(Feedback[41]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U2 ( .A1(PermutationOutput[40]), 
        .A2(PermutationOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_1_U1 ( .A1(PermutationOutput[40]), .A2(
        PermutationOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_10_LFInst_2_U2 ( .B1(PermutationOutput[43]), 
        .B2(PermutationOutput[40]), .A(SubCellInst_LFInst_10_LFInst_2_n1), 
        .ZN(Feedback[42]) );
  OAI221_X1 SubCellInst_LFInst_10_LFInst_2_U1 ( .B1(PermutationOutput[42]), 
        .B2(PermutationOutput[43]), .C1(PermutationOutput[42]), .C2(
        PermutationOutput[40]), .A(PermutationOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_10_LFInst_3_U1 ( .A1(PermutationOutput[41]), 
        .A2(PermutationOutput[43]), .B1(PermutationOutput[41]), .B2(
        PermutationOutput[40]), .C1(PermutationOutput[43]), .C2(
        PermutationOutput[42]), .ZN(Feedback[43]) );
  AOI21_X1 SubCellInst_LFInst_11_LFInst_0_U2 ( .B1(PermutationOutput[47]), 
        .B2(PermutationOutput[46]), .A(SubCellInst_LFInst_11_LFInst_0_n1), 
        .ZN(Feedback[44]) );
  AOI221_X1 SubCellInst_LFInst_11_LFInst_0_U1 ( .B1(PermutationOutput[46]), 
        .B2(PermutationOutput[44]), .C1(PermutationOutput[47]), .C2(
        PermutationOutput[44]), .A(PermutationOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_11_LFInst_1_U3 ( .B1(PermutationOutput[47]), 
        .B2(SubCellInst_LFInst_11_LFInst_1_n2), .A(
        SubCellInst_LFInst_11_LFInst_1_n1), .ZN(Feedback[45]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U2 ( .A1(PermutationOutput[44]), 
        .A2(PermutationOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_1_U1 ( .A1(PermutationOutput[44]), .A2(
        PermutationOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_11_LFInst_2_U2 ( .B1(PermutationOutput[47]), 
        .B2(PermutationOutput[44]), .A(SubCellInst_LFInst_11_LFInst_2_n1), 
        .ZN(Feedback[46]) );
  OAI221_X1 SubCellInst_LFInst_11_LFInst_2_U1 ( .B1(PermutationOutput[46]), 
        .B2(PermutationOutput[47]), .C1(PermutationOutput[46]), .C2(
        PermutationOutput[44]), .A(PermutationOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_11_LFInst_3_U1 ( .A1(PermutationOutput[45]), 
        .A2(PermutationOutput[47]), .B1(PermutationOutput[45]), .B2(
        PermutationOutput[44]), .C1(PermutationOutput[47]), .C2(
        PermutationOutput[46]), .ZN(Feedback[47]) );
  AOI21_X1 SubCellInst_LFInst_12_LFInst_0_U2 ( .B1(PermutationOutput[51]), 
        .B2(PermutationOutput[50]), .A(SubCellInst_LFInst_12_LFInst_0_n1), 
        .ZN(Feedback[48]) );
  AOI221_X1 SubCellInst_LFInst_12_LFInst_0_U1 ( .B1(PermutationOutput[50]), 
        .B2(PermutationOutput[48]), .C1(PermutationOutput[51]), .C2(
        PermutationOutput[48]), .A(PermutationOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_12_LFInst_1_U3 ( .B1(PermutationOutput[51]), 
        .B2(SubCellInst_LFInst_12_LFInst_1_n2), .A(
        SubCellInst_LFInst_12_LFInst_1_n1), .ZN(Feedback[49]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U2 ( .A1(PermutationOutput[48]), 
        .A2(PermutationOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_1_U1 ( .A1(PermutationOutput[48]), .A2(
        PermutationOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_12_LFInst_2_U2 ( .B1(PermutationOutput[51]), 
        .B2(PermutationOutput[48]), .A(SubCellInst_LFInst_12_LFInst_2_n1), 
        .ZN(Feedback[50]) );
  OAI221_X1 SubCellInst_LFInst_12_LFInst_2_U1 ( .B1(PermutationOutput[50]), 
        .B2(PermutationOutput[51]), .C1(PermutationOutput[50]), .C2(
        PermutationOutput[48]), .A(PermutationOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_12_LFInst_3_U1 ( .A1(PermutationOutput[49]), 
        .A2(PermutationOutput[51]), .B1(PermutationOutput[49]), .B2(
        PermutationOutput[48]), .C1(PermutationOutput[51]), .C2(
        PermutationOutput[50]), .ZN(Feedback[51]) );
  AOI21_X1 SubCellInst_LFInst_13_LFInst_0_U2 ( .B1(PermutationOutput[55]), 
        .B2(PermutationOutput[54]), .A(SubCellInst_LFInst_13_LFInst_0_n1), 
        .ZN(Feedback[52]) );
  AOI221_X1 SubCellInst_LFInst_13_LFInst_0_U1 ( .B1(PermutationOutput[54]), 
        .B2(PermutationOutput[52]), .C1(PermutationOutput[55]), .C2(
        PermutationOutput[52]), .A(PermutationOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_13_LFInst_1_U3 ( .B1(PermutationOutput[55]), 
        .B2(SubCellInst_LFInst_13_LFInst_1_n2), .A(
        SubCellInst_LFInst_13_LFInst_1_n1), .ZN(Feedback[53]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U2 ( .A1(PermutationOutput[52]), 
        .A2(PermutationOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_1_U1 ( .A1(PermutationOutput[52]), .A2(
        PermutationOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_13_LFInst_2_U2 ( .B1(PermutationOutput[55]), 
        .B2(PermutationOutput[52]), .A(SubCellInst_LFInst_13_LFInst_2_n1), 
        .ZN(Feedback[54]) );
  OAI221_X1 SubCellInst_LFInst_13_LFInst_2_U1 ( .B1(PermutationOutput[54]), 
        .B2(PermutationOutput[55]), .C1(PermutationOutput[54]), .C2(
        PermutationOutput[52]), .A(PermutationOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_13_LFInst_3_U1 ( .A1(PermutationOutput[53]), 
        .A2(PermutationOutput[55]), .B1(PermutationOutput[53]), .B2(
        PermutationOutput[52]), .C1(PermutationOutput[55]), .C2(
        PermutationOutput[54]), .ZN(Feedback[55]) );
  AOI21_X1 SubCellInst_LFInst_14_LFInst_0_U2 ( .B1(PermutationOutput[59]), 
        .B2(PermutationOutput[58]), .A(SubCellInst_LFInst_14_LFInst_0_n1), 
        .ZN(Feedback[56]) );
  AOI221_X1 SubCellInst_LFInst_14_LFInst_0_U1 ( .B1(PermutationOutput[58]), 
        .B2(PermutationOutput[56]), .C1(PermutationOutput[59]), .C2(
        PermutationOutput[56]), .A(PermutationOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_14_LFInst_1_U3 ( .B1(PermutationOutput[59]), 
        .B2(SubCellInst_LFInst_14_LFInst_1_n2), .A(
        SubCellInst_LFInst_14_LFInst_1_n1), .ZN(Feedback[57]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U2 ( .A1(PermutationOutput[56]), 
        .A2(PermutationOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_1_U1 ( .A1(PermutationOutput[56]), .A2(
        PermutationOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_14_LFInst_2_U2 ( .B1(PermutationOutput[59]), 
        .B2(PermutationOutput[56]), .A(SubCellInst_LFInst_14_LFInst_2_n1), 
        .ZN(Feedback[58]) );
  OAI221_X1 SubCellInst_LFInst_14_LFInst_2_U1 ( .B1(PermutationOutput[58]), 
        .B2(PermutationOutput[59]), .C1(PermutationOutput[58]), .C2(
        PermutationOutput[56]), .A(PermutationOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_14_LFInst_3_U1 ( .A1(PermutationOutput[57]), 
        .A2(PermutationOutput[59]), .B1(PermutationOutput[57]), .B2(
        PermutationOutput[56]), .C1(PermutationOutput[59]), .C2(
        PermutationOutput[58]), .ZN(Feedback[59]) );
  AOI21_X1 SubCellInst_LFInst_15_LFInst_0_U2 ( .B1(PermutationOutput[63]), 
        .B2(PermutationOutput[62]), .A(SubCellInst_LFInst_15_LFInst_0_n1), 
        .ZN(Feedback[60]) );
  AOI221_X1 SubCellInst_LFInst_15_LFInst_0_U1 ( .B1(PermutationOutput[62]), 
        .B2(PermutationOutput[60]), .C1(PermutationOutput[63]), .C2(
        PermutationOutput[60]), .A(PermutationOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n1) );
  OAI21_X1 SubCellInst_LFInst_15_LFInst_1_U3 ( .B1(PermutationOutput[63]), 
        .B2(SubCellInst_LFInst_15_LFInst_1_n2), .A(
        SubCellInst_LFInst_15_LFInst_1_n1), .ZN(Feedback[61]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U2 ( .A1(PermutationOutput[60]), 
        .A2(PermutationOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_1_n1) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_1_U1 ( .A1(PermutationOutput[60]), .A2(
        PermutationOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_1_n2) );
  OAI21_X1 SubCellInst_LFInst_15_LFInst_2_U2 ( .B1(PermutationOutput[63]), 
        .B2(PermutationOutput[60]), .A(SubCellInst_LFInst_15_LFInst_2_n1), 
        .ZN(Feedback[62]) );
  OAI221_X1 SubCellInst_LFInst_15_LFInst_2_U1 ( .B1(PermutationOutput[62]), 
        .B2(PermutationOutput[63]), .C1(PermutationOutput[62]), .C2(
        PermutationOutput[60]), .A(PermutationOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n1) );
  AOI222_X1 SubCellInst_LFInst_15_LFInst_3_U1 ( .A1(PermutationOutput[61]), 
        .A2(PermutationOutput[63]), .B1(PermutationOutput[61]), .B2(
        PermutationOutput[60]), .C1(PermutationOutput[63]), .C2(
        PermutationOutput[62]), .ZN(Feedback[63]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_0_n1), .B(Input[2]), .ZN(
        Red_Input[0]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U1 ( .A(Input[0]), .B(Input[1]), 
        .ZN(Red_PlaintextInst_LFInst_0_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_1_n1), .B(Input[3]), .ZN(
        Red_Input[1]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_1_U1 ( .A(Input[0]), .B(Input[1]), 
        .ZN(Red_PlaintextInst_LFInst_0_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_2_n1), .B(Input[3]), .ZN(
        Red_Input[2]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_2_U1 ( .A(Input[1]), .B(Input[2]), 
        .ZN(Red_PlaintextInst_LFInst_0_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_0_n1), .B(Input[6]), .ZN(
        Red_Input[3]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U1 ( .A(Input[4]), .B(Input[5]), 
        .ZN(Red_PlaintextInst_LFInst_1_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_1_n1), .B(Input[7]), .ZN(
        Red_Input[4]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_1_U1 ( .A(Input[4]), .B(Input[5]), 
        .ZN(Red_PlaintextInst_LFInst_1_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_2_n1), .B(Input[7]), .ZN(
        Red_Input[5]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_2_U1 ( .A(Input[5]), .B(Input[6]), 
        .ZN(Red_PlaintextInst_LFInst_1_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_0_n1), .B(Input[10]), .ZN(
        Red_Input[6]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U1 ( .A(Input[8]), .B(Input[9]), 
        .ZN(Red_PlaintextInst_LFInst_2_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_1_n1), .B(Input[11]), .ZN(
        Red_Input[7]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_1_U1 ( .A(Input[8]), .B(Input[9]), 
        .ZN(Red_PlaintextInst_LFInst_2_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_2_n1), .B(Input[11]), .ZN(
        Red_Input[8]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_2_U1 ( .A(Input[9]), .B(Input[10]), .ZN(Red_PlaintextInst_LFInst_2_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_0_n1), .B(Input[14]), .ZN(
        Red_Input[9]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U1 ( .A(Input[12]), .B(
        Input[13]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_1_n1), .B(Input[15]), .ZN(
        Red_Input[10]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_1_U1 ( .A(Input[12]), .B(
        Input[13]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_2_n1), .B(Input[15]), .ZN(
        Red_Input[11]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_2_U1 ( .A(Input[13]), .B(
        Input[14]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_0_n1), .B(Input[18]), .ZN(
        Red_Input[12]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U1 ( .A(Input[16]), .B(
        Input[17]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_1_n1), .B(Input[19]), .ZN(
        Red_Input[13]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_1_U1 ( .A(Input[16]), .B(
        Input[17]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_2_n1), .B(Input[19]), .ZN(
        Red_Input[14]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_2_U1 ( .A(Input[17]), .B(
        Input[18]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_0_n1), .B(Input[22]), .ZN(
        Red_Input[15]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U1 ( .A(Input[20]), .B(
        Input[21]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_1_n1), .B(Input[23]), .ZN(
        Red_Input[16]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_1_U1 ( .A(Input[20]), .B(
        Input[21]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_2_n1), .B(Input[23]), .ZN(
        Red_Input[17]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_2_U1 ( .A(Input[21]), .B(
        Input[22]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_0_n1), .B(Input[26]), .ZN(
        Red_Input[18]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U1 ( .A(Input[24]), .B(
        Input[25]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_1_n1), .B(Input[27]), .ZN(
        Red_Input[19]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_1_U1 ( .A(Input[24]), .B(
        Input[25]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_2_n1), .B(Input[27]), .ZN(
        Red_Input[20]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_2_U1 ( .A(Input[25]), .B(
        Input[26]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_0_n1), .B(Input[30]), .ZN(
        Red_Input[21]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U1 ( .A(Input[28]), .B(
        Input[29]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_1_n1), .B(Input[31]), .ZN(
        Red_Input[22]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_1_U1 ( .A(Input[28]), .B(
        Input[29]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_2_n1), .B(Input[31]), .ZN(
        Red_Input[23]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_2_U1 ( .A(Input[29]), .B(
        Input[30]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_0_n1), .B(Input[34]), .ZN(
        Red_Input[24]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U1 ( .A(Input[32]), .B(
        Input[33]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_1_n1), .B(Input[35]), .ZN(
        Red_Input[25]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_1_U1 ( .A(Input[32]), .B(
        Input[33]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_2_n1), .B(Input[35]), .ZN(
        Red_Input[26]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_2_U1 ( .A(Input[33]), .B(
        Input[34]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_0_n1), .B(Input[38]), .ZN(
        Red_Input[27]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U1 ( .A(Input[36]), .B(
        Input[37]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_1_n1), .B(Input[39]), .ZN(
        Red_Input[28]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_1_U1 ( .A(Input[36]), .B(
        Input[37]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_2_n1), .B(Input[39]), .ZN(
        Red_Input[29]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_2_U1 ( .A(Input[37]), .B(
        Input[38]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_0_n1), .B(Input[42]), .ZN(
        Red_Input[30]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U1 ( .A(Input[40]), .B(
        Input[41]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_1_n1), .B(Input[43]), .ZN(
        Red_Input[31]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_1_U1 ( .A(Input[40]), .B(
        Input[41]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_2_n1), .B(Input[43]), .ZN(
        Red_Input[32]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_2_U1 ( .A(Input[41]), .B(
        Input[42]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_0_n1), .B(Input[46]), .ZN(
        Red_Input[33]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U1 ( .A(Input[44]), .B(
        Input[45]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_1_n1), .B(Input[47]), .ZN(
        Red_Input[34]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_1_U1 ( .A(Input[44]), .B(
        Input[45]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_2_n1), .B(Input[47]), .ZN(
        Red_Input[35]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_2_U1 ( .A(Input[45]), .B(
        Input[46]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_0_n1), .B(Input[50]), .ZN(
        Red_Input[36]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U1 ( .A(Input[48]), .B(
        Input[49]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_1_n1), .B(Input[51]), .ZN(
        Red_Input[37]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_1_U1 ( .A(Input[48]), .B(
        Input[49]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_2_n1), .B(Input[51]), .ZN(
        Red_Input[38]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_2_U1 ( .A(Input[49]), .B(
        Input[50]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_0_n1), .B(Input[54]), .ZN(
        Red_Input[39]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U1 ( .A(Input[52]), .B(
        Input[53]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_1_n1), .B(Input[55]), .ZN(
        Red_Input[40]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_1_U1 ( .A(Input[52]), .B(
        Input[53]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_2_n1), .B(Input[55]), .ZN(
        Red_Input[41]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_2_U1 ( .A(Input[53]), .B(
        Input[54]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_0_n1), .B(Input[58]), .ZN(
        Red_Input[42]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U1 ( .A(Input[56]), .B(
        Input[57]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_1_n1), .B(Input[59]), .ZN(
        Red_Input[43]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_1_U1 ( .A(Input[56]), .B(
        Input[57]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_2_n1), .B(Input[59]), .ZN(
        Red_Input[44]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_2_U1 ( .A(Input[57]), .B(
        Input[58]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_2_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_0_n1), .B(Input[62]), .ZN(
        Red_Input[45]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U1 ( .A(Input[60]), .B(
        Input[61]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_0_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_1_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_1_n1), .B(Input[63]), .ZN(
        Red_Input[46]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_1_U1 ( .A(Input[60]), .B(
        Input[61]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_1_n1) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_2_U2 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_2_n1), .B(Input[63]), .ZN(
        Red_Input[47]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_2_U1 ( .A(Input[61]), .B(
        Input[62]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_2_n1) );
  MUX2_X1 Red_InputMUX_MUXInst_0_U1 ( .A(Red_Feedback[0]), .B(Red_Input[0]), 
        .S(rst), .Z(Red_MCOutput[0]) );
  MUX2_X1 Red_InputMUX_MUXInst_1_U1 ( .A(Red_Feedback[1]), .B(Red_Input[1]), 
        .S(rst), .Z(Red_MCOutput[1]) );
  MUX2_X1 Red_InputMUX_MUXInst_2_U1 ( .A(Red_Feedback[2]), .B(Red_Input[2]), 
        .S(rst), .Z(Red_MCOutput[2]) );
  MUX2_X1 Red_InputMUX_MUXInst_3_U1 ( .A(Red_Feedback[3]), .B(Red_Input[3]), 
        .S(rst), .Z(Red_MCOutput[3]) );
  MUX2_X1 Red_InputMUX_MUXInst_4_U1 ( .A(Red_Feedback[4]), .B(Red_Input[4]), 
        .S(rst), .Z(Red_MCOutput[4]) );
  MUX2_X1 Red_InputMUX_MUXInst_5_U1 ( .A(Red_Feedback[5]), .B(Red_Input[5]), 
        .S(rst), .Z(Red_MCOutput[5]) );
  MUX2_X1 Red_InputMUX_MUXInst_6_U1 ( .A(Red_Feedback[6]), .B(Red_Input[6]), 
        .S(rst), .Z(Red_MCOutput[6]) );
  MUX2_X1 Red_InputMUX_MUXInst_7_U1 ( .A(Red_Feedback[7]), .B(Red_Input[7]), 
        .S(rst), .Z(Red_MCOutput[7]) );
  MUX2_X1 Red_InputMUX_MUXInst_8_U1 ( .A(Red_Feedback[8]), .B(Red_Input[8]), 
        .S(rst), .Z(Red_MCOutput[8]) );
  MUX2_X1 Red_InputMUX_MUXInst_9_U1 ( .A(Red_Feedback[9]), .B(Red_Input[9]), 
        .S(rst), .Z(Red_MCOutput[9]) );
  MUX2_X1 Red_InputMUX_MUXInst_10_U1 ( .A(Red_Feedback[10]), .B(Red_Input[10]), 
        .S(rst), .Z(Red_MCOutput[10]) );
  MUX2_X1 Red_InputMUX_MUXInst_11_U1 ( .A(Red_Feedback[11]), .B(Red_Input[11]), 
        .S(rst), .Z(Red_MCOutput[11]) );
  MUX2_X1 Red_InputMUX_MUXInst_12_U1 ( .A(Red_Feedback[12]), .B(Red_Input[12]), 
        .S(rst), .Z(Red_MCOutput[12]) );
  MUX2_X1 Red_InputMUX_MUXInst_13_U1 ( .A(Red_Feedback[13]), .B(Red_Input[13]), 
        .S(rst), .Z(Red_MCOutput[13]) );
  MUX2_X1 Red_InputMUX_MUXInst_14_U1 ( .A(Red_Feedback[14]), .B(Red_Input[14]), 
        .S(rst), .Z(Red_MCOutput[14]) );
  MUX2_X1 Red_InputMUX_MUXInst_15_U1 ( .A(Red_Feedback[15]), .B(Red_Input[15]), 
        .S(rst), .Z(Red_MCOutput[15]) );
  MUX2_X1 Red_InputMUX_MUXInst_16_U1 ( .A(Red_Feedback[16]), .B(Red_Input[16]), 
        .S(rst), .Z(Red_MCOutput[16]) );
  MUX2_X1 Red_InputMUX_MUXInst_17_U1 ( .A(Red_Feedback[17]), .B(Red_Input[17]), 
        .S(rst), .Z(Red_MCOutput[17]) );
  MUX2_X1 Red_InputMUX_MUXInst_18_U1 ( .A(Red_Feedback[18]), .B(Red_Input[18]), 
        .S(rst), .Z(Red_MCOutput[18]) );
  MUX2_X1 Red_InputMUX_MUXInst_19_U1 ( .A(Red_Feedback[19]), .B(Red_Input[19]), 
        .S(rst), .Z(Red_MCOutput[19]) );
  MUX2_X1 Red_InputMUX_MUXInst_20_U1 ( .A(Red_Feedback[20]), .B(Red_Input[20]), 
        .S(rst), .Z(Red_MCOutput[20]) );
  MUX2_X1 Red_InputMUX_MUXInst_21_U1 ( .A(Red_Feedback[21]), .B(Red_Input[21]), 
        .S(rst), .Z(Red_MCOutput[21]) );
  MUX2_X1 Red_InputMUX_MUXInst_22_U1 ( .A(Red_Feedback[22]), .B(Red_Input[22]), 
        .S(rst), .Z(Red_MCOutput[22]) );
  MUX2_X1 Red_InputMUX_MUXInst_23_U1 ( .A(Red_Feedback[23]), .B(Red_Input[23]), 
        .S(rst), .Z(Red_MCOutput[23]) );
  MUX2_X1 Red_InputMUX_MUXInst_24_U1 ( .A(Red_Feedback[24]), .B(Red_Input[24]), 
        .S(rst), .Z(Red_MCInput[24]) );
  MUX2_X1 Red_InputMUX_MUXInst_25_U1 ( .A(Red_Feedback[25]), .B(Red_Input[25]), 
        .S(rst), .Z(Red_MCInput[25]) );
  MUX2_X1 Red_InputMUX_MUXInst_26_U1 ( .A(Red_Feedback[26]), .B(Red_Input[26]), 
        .S(rst), .Z(Red_MCInput[26]) );
  MUX2_X1 Red_InputMUX_MUXInst_27_U1 ( .A(Red_Feedback[27]), .B(Red_Input[27]), 
        .S(rst), .Z(Red_MCInput[27]) );
  MUX2_X1 Red_InputMUX_MUXInst_28_U1 ( .A(Red_Feedback[28]), .B(Red_Input[28]), 
        .S(rst), .Z(Red_MCInput[28]) );
  MUX2_X1 Red_InputMUX_MUXInst_29_U1 ( .A(Red_Feedback[29]), .B(Red_Input[29]), 
        .S(rst), .Z(Red_MCInput[29]) );
  MUX2_X1 Red_InputMUX_MUXInst_30_U1 ( .A(Red_Feedback[30]), .B(Red_Input[30]), 
        .S(rst), .Z(Red_MCInput[30]) );
  MUX2_X1 Red_InputMUX_MUXInst_31_U1 ( .A(Red_Feedback[31]), .B(Red_Input[31]), 
        .S(rst), .Z(Red_MCInput[31]) );
  MUX2_X1 Red_InputMUX_MUXInst_32_U1 ( .A(Red_Feedback[32]), .B(Red_Input[32]), 
        .S(rst), .Z(Red_MCInput[32]) );
  MUX2_X1 Red_InputMUX_MUXInst_33_U1 ( .A(Red_Feedback[33]), .B(Red_Input[33]), 
        .S(rst), .Z(Red_MCInput[33]) );
  MUX2_X1 Red_InputMUX_MUXInst_34_U1 ( .A(Red_Feedback[34]), .B(Red_Input[34]), 
        .S(rst), .Z(Red_MCInput[34]) );
  MUX2_X1 Red_InputMUX_MUXInst_35_U1 ( .A(Red_Feedback[35]), .B(Red_Input[35]), 
        .S(rst), .Z(Red_MCInput[35]) );
  MUX2_X1 Red_InputMUX_MUXInst_36_U1 ( .A(Red_Feedback[36]), .B(Red_Input[36]), 
        .S(rst), .Z(Red_MCInput[36]) );
  MUX2_X1 Red_InputMUX_MUXInst_37_U1 ( .A(Red_Feedback[37]), .B(Red_Input[37]), 
        .S(rst), .Z(Red_MCInput[37]) );
  MUX2_X1 Red_InputMUX_MUXInst_38_U1 ( .A(Red_Feedback[38]), .B(Red_Input[38]), 
        .S(rst), .Z(Red_MCInput[38]) );
  MUX2_X1 Red_InputMUX_MUXInst_39_U1 ( .A(Red_Feedback[39]), .B(Red_Input[39]), 
        .S(rst), .Z(Red_MCInput[39]) );
  MUX2_X1 Red_InputMUX_MUXInst_40_U1 ( .A(Red_Feedback[40]), .B(Red_Input[40]), 
        .S(rst), .Z(Red_MCInput[40]) );
  MUX2_X1 Red_InputMUX_MUXInst_41_U1 ( .A(Red_Feedback[41]), .B(Red_Input[41]), 
        .S(rst), .Z(Red_MCInput[41]) );
  MUX2_X1 Red_InputMUX_MUXInst_42_U1 ( .A(Red_Feedback[42]), .B(Red_Input[42]), 
        .S(rst), .Z(Red_MCInput[42]) );
  MUX2_X1 Red_InputMUX_MUXInst_43_U1 ( .A(Red_Feedback[43]), .B(Red_Input[43]), 
        .S(rst), .Z(Red_MCInput[43]) );
  MUX2_X1 Red_InputMUX_MUXInst_44_U1 ( .A(Red_Feedback[44]), .B(Red_Input[44]), 
        .S(rst), .Z(Red_MCInput[44]) );
  MUX2_X1 Red_InputMUX_MUXInst_45_U1 ( .A(Red_Feedback[45]), .B(Red_Input[45]), 
        .S(rst), .Z(Red_MCInput[45]) );
  MUX2_X1 Red_InputMUX_MUXInst_46_U1 ( .A(Red_Feedback[46]), .B(Red_Input[46]), 
        .S(rst), .Z(Red_MCInput[46]) );
  MUX2_X1 Red_InputMUX_MUXInst_47_U1 ( .A(Red_Feedback[47]), .B(Red_Input[47]), 
        .S(rst), .Z(Red_MCInput[47]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_0_U3 ( .A(Red_MCInst_XOR_r0_Inst_0_n2), .B(
        Red_MCInst_XOR_r0_Inst_0_n1), .ZN(Red_MCOutput[36]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_0_U2 ( .A(Red_MCOutput[12]), .B(
        Red_MCOutput[0]), .ZN(Red_MCInst_XOR_r0_Inst_0_n1) );
  XOR2_X1 Red_MCInst_XOR_r0_Inst_0_U1 ( .A(1'b0), .B(Red_MCInput[36]), .Z(
        Red_MCInst_XOR_r0_Inst_0_n2) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_0_U2 ( .A(Red_MCInst_XOR_r1_Inst_0_n1), .B(
        Red_MCOutput[0]), .ZN(Red_MCOutput[24]) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_0_U1 ( .A(1'b0), .B(Red_MCInput[24]), .ZN(
        Red_MCInst_XOR_r1_Inst_0_n1) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_1_U3 ( .A(Red_MCInst_XOR_r0_Inst_1_n2), .B(
        Red_MCInst_XOR_r0_Inst_1_n1), .ZN(Red_MCOutput[37]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_1_U2 ( .A(Red_MCOutput[13]), .B(
        Red_MCOutput[1]), .ZN(Red_MCInst_XOR_r0_Inst_1_n1) );
  XOR2_X1 Red_MCInst_XOR_r0_Inst_1_U1 ( .A(1'b0), .B(Red_MCInput[37]), .Z(
        Red_MCInst_XOR_r0_Inst_1_n2) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_1_U2 ( .A(Red_MCInst_XOR_r1_Inst_1_n1), .B(
        Red_MCOutput[1]), .ZN(Red_MCOutput[25]) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_1_U1 ( .A(1'b0), .B(Red_MCInput[25]), .ZN(
        Red_MCInst_XOR_r1_Inst_1_n1) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_2_U3 ( .A(Red_MCInst_XOR_r0_Inst_2_n2), .B(
        Red_MCInst_XOR_r0_Inst_2_n1), .ZN(Red_MCOutput[38]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_2_U2 ( .A(Red_MCOutput[14]), .B(
        Red_MCOutput[2]), .ZN(Red_MCInst_XOR_r0_Inst_2_n1) );
  XOR2_X1 Red_MCInst_XOR_r0_Inst_2_U1 ( .A(1'b0), .B(Red_MCInput[38]), .Z(
        Red_MCInst_XOR_r0_Inst_2_n2) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_2_U2 ( .A(Red_MCInst_XOR_r1_Inst_2_n1), .B(
        Red_MCOutput[2]), .ZN(Red_MCOutput[26]) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_2_U1 ( .A(1'b0), .B(Red_MCInput[26]), .ZN(
        Red_MCInst_XOR_r1_Inst_2_n1) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_3_U3 ( .A(Red_MCInst_XOR_r0_Inst_3_n2), .B(
        Red_MCInst_XOR_r0_Inst_3_n1), .ZN(Red_MCOutput[39]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_3_U2 ( .A(Red_MCOutput[15]), .B(
        Red_MCOutput[3]), .ZN(Red_MCInst_XOR_r0_Inst_3_n1) );
  XOR2_X1 Red_MCInst_XOR_r0_Inst_3_U1 ( .A(1'b0), .B(Red_MCInput[39]), .Z(
        Red_MCInst_XOR_r0_Inst_3_n2) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_3_U2 ( .A(Red_MCInst_XOR_r1_Inst_3_n1), .B(
        Red_MCOutput[3]), .ZN(Red_MCOutput[27]) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_3_U1 ( .A(1'b0), .B(Red_MCInput[27]), .ZN(
        Red_MCInst_XOR_r1_Inst_3_n1) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_4_U3 ( .A(Red_MCInst_XOR_r0_Inst_4_n2), .B(
        Red_MCInst_XOR_r0_Inst_4_n1), .ZN(Red_MCOutput[40]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_4_U2 ( .A(Red_MCOutput[16]), .B(
        Red_MCOutput[4]), .ZN(Red_MCInst_XOR_r0_Inst_4_n1) );
  XOR2_X1 Red_MCInst_XOR_r0_Inst_4_U1 ( .A(1'b0), .B(Red_MCInput[40]), .Z(
        Red_MCInst_XOR_r0_Inst_4_n2) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_4_U2 ( .A(Red_MCInst_XOR_r1_Inst_4_n1), .B(
        Red_MCOutput[4]), .ZN(Red_MCOutput[28]) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_4_U1 ( .A(1'b0), .B(Red_MCInput[28]), .ZN(
        Red_MCInst_XOR_r1_Inst_4_n1) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_5_U3 ( .A(Red_MCInst_XOR_r0_Inst_5_n2), .B(
        Red_MCInst_XOR_r0_Inst_5_n1), .ZN(Red_MCOutput[41]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_5_U2 ( .A(Red_MCOutput[17]), .B(
        Red_MCOutput[5]), .ZN(Red_MCInst_XOR_r0_Inst_5_n1) );
  XOR2_X1 Red_MCInst_XOR_r0_Inst_5_U1 ( .A(1'b0), .B(Red_MCInput[41]), .Z(
        Red_MCInst_XOR_r0_Inst_5_n2) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_5_U2 ( .A(Red_MCInst_XOR_r1_Inst_5_n1), .B(
        Red_MCOutput[5]), .ZN(Red_MCOutput[29]) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_5_U1 ( .A(1'b0), .B(Red_MCInput[29]), .ZN(
        Red_MCInst_XOR_r1_Inst_5_n1) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_6_U3 ( .A(Red_MCInst_XOR_r0_Inst_6_n2), .B(
        Red_MCInst_XOR_r0_Inst_6_n1), .ZN(Red_MCOutput[42]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_6_U2 ( .A(Red_MCOutput[18]), .B(
        Red_MCOutput[6]), .ZN(Red_MCInst_XOR_r0_Inst_6_n1) );
  XOR2_X1 Red_MCInst_XOR_r0_Inst_6_U1 ( .A(1'b0), .B(Red_MCInput[42]), .Z(
        Red_MCInst_XOR_r0_Inst_6_n2) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_6_U2 ( .A(Red_MCInst_XOR_r1_Inst_6_n1), .B(
        Red_MCOutput[6]), .ZN(Red_MCOutput[30]) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_6_U1 ( .A(1'b0), .B(Red_MCInput[30]), .ZN(
        Red_MCInst_XOR_r1_Inst_6_n1) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_7_U3 ( .A(Red_MCInst_XOR_r0_Inst_7_n2), .B(
        Red_MCInst_XOR_r0_Inst_7_n1), .ZN(Red_MCOutput[43]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_7_U2 ( .A(Red_MCOutput[19]), .B(
        Red_MCOutput[7]), .ZN(Red_MCInst_XOR_r0_Inst_7_n1) );
  XOR2_X1 Red_MCInst_XOR_r0_Inst_7_U1 ( .A(1'b0), .B(Red_MCInput[43]), .Z(
        Red_MCInst_XOR_r0_Inst_7_n2) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_7_U2 ( .A(Red_MCInst_XOR_r1_Inst_7_n1), .B(
        Red_MCOutput[7]), .ZN(Red_MCOutput[31]) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_7_U1 ( .A(1'b0), .B(Red_MCInput[31]), .ZN(
        Red_MCInst_XOR_r1_Inst_7_n1) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_8_U3 ( .A(Red_MCInst_XOR_r0_Inst_8_n2), .B(
        Red_MCInst_XOR_r0_Inst_8_n1), .ZN(Red_MCOutput[44]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_8_U2 ( .A(Red_MCOutput[20]), .B(
        Red_MCOutput[8]), .ZN(Red_MCInst_XOR_r0_Inst_8_n1) );
  XOR2_X1 Red_MCInst_XOR_r0_Inst_8_U1 ( .A(1'b0), .B(Red_MCInput[44]), .Z(
        Red_MCInst_XOR_r0_Inst_8_n2) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_8_U2 ( .A(Red_MCInst_XOR_r1_Inst_8_n1), .B(
        Red_MCOutput[8]), .ZN(Red_MCOutput[32]) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_8_U1 ( .A(1'b0), .B(Red_MCInput[32]), .ZN(
        Red_MCInst_XOR_r1_Inst_8_n1) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_9_U3 ( .A(Red_MCInst_XOR_r0_Inst_9_n2), .B(
        Red_MCInst_XOR_r0_Inst_9_n1), .ZN(Red_MCOutput[45]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_9_U2 ( .A(Red_MCOutput[21]), .B(
        Red_MCOutput[9]), .ZN(Red_MCInst_XOR_r0_Inst_9_n1) );
  XOR2_X1 Red_MCInst_XOR_r0_Inst_9_U1 ( .A(1'b0), .B(Red_MCInput[45]), .Z(
        Red_MCInst_XOR_r0_Inst_9_n2) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_9_U2 ( .A(Red_MCInst_XOR_r1_Inst_9_n1), .B(
        Red_MCOutput[9]), .ZN(Red_MCOutput[33]) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_9_U1 ( .A(1'b0), .B(Red_MCInput[33]), .ZN(
        Red_MCInst_XOR_r1_Inst_9_n1) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_10_U3 ( .A(Red_MCInst_XOR_r0_Inst_10_n2), 
        .B(Red_MCInst_XOR_r0_Inst_10_n1), .ZN(Red_MCOutput[46]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_10_U2 ( .A(Red_MCOutput[22]), .B(
        Red_MCOutput[10]), .ZN(Red_MCInst_XOR_r0_Inst_10_n1) );
  XOR2_X1 Red_MCInst_XOR_r0_Inst_10_U1 ( .A(1'b0), .B(Red_MCInput[46]), .Z(
        Red_MCInst_XOR_r0_Inst_10_n2) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_10_U2 ( .A(Red_MCInst_XOR_r1_Inst_10_n1), 
        .B(Red_MCOutput[10]), .ZN(Red_MCOutput[34]) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_10_U1 ( .A(1'b0), .B(Red_MCInput[34]), .ZN(
        Red_MCInst_XOR_r1_Inst_10_n1) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_11_U3 ( .A(Red_MCInst_XOR_r0_Inst_11_n2), 
        .B(Red_MCInst_XOR_r0_Inst_11_n1), .ZN(Red_MCOutput[47]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_11_U2 ( .A(Red_MCOutput[23]), .B(
        Red_MCOutput[11]), .ZN(Red_MCInst_XOR_r0_Inst_11_n1) );
  XOR2_X1 Red_MCInst_XOR_r0_Inst_11_U1 ( .A(1'b0), .B(Red_MCInput[47]), .Z(
        Red_MCInst_XOR_r0_Inst_11_n2) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_11_U2 ( .A(Red_MCInst_XOR_r1_Inst_11_n1), 
        .B(Red_MCOutput[11]), .ZN(Red_MCOutput[35]) );
  XNOR2_X1 Red_MCInst_XOR_r1_Inst_11_U1 ( .A(1'b0), .B(Red_MCInput[35]), .ZN(
        Red_MCInst_XOR_r1_Inst_11_n1) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_0_0_U2 ( .A(Red_AddKeyXOR1_XORInst_0_0_n1), 
        .B(Red_SelectedKey[36]), .ZN(Red_final[36]) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_0_0_U1 ( .A(1'b0), .B(Red_MCOutput[36]), 
        .ZN(Red_AddKeyXOR1_XORInst_0_0_n1) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_0_1_U2 ( .A(Red_AddKeyXOR1_XORInst_0_1_n1), 
        .B(Red_SelectedKey[37]), .ZN(Red_final[37]) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_0_1_U1 ( .A(1'b0), .B(Red_MCOutput[37]), 
        .ZN(Red_AddKeyXOR1_XORInst_0_1_n1) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_0_2_U2 ( .A(Red_AddKeyXOR1_XORInst_0_2_n1), 
        .B(Red_SelectedKey[38]), .ZN(Red_final[38]) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_0_2_U1 ( .A(1'b0), .B(Red_MCOutput[38]), 
        .ZN(Red_AddKeyXOR1_XORInst_0_2_n1) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_1_0_U2 ( .A(Red_AddKeyXOR1_XORInst_1_0_n1), 
        .B(Red_SelectedKey[39]), .ZN(Red_final[39]) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_1_0_U1 ( .A(1'b0), .B(Red_MCOutput[39]), 
        .ZN(Red_AddKeyXOR1_XORInst_1_0_n1) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_1_1_U2 ( .A(Red_AddKeyXOR1_XORInst_1_1_n1), 
        .B(Red_SelectedKey[40]), .ZN(Red_final[40]) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_1_1_U1 ( .A(1'b0), .B(Red_MCOutput[40]), 
        .ZN(Red_AddKeyXOR1_XORInst_1_1_n1) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_1_2_U2 ( .A(Red_AddKeyXOR1_XORInst_1_2_n1), 
        .B(Red_SelectedKey[41]), .ZN(Red_final[41]) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_1_2_U1 ( .A(1'b0), .B(Red_MCOutput[41]), 
        .ZN(Red_AddKeyXOR1_XORInst_1_2_n1) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_2_0_U2 ( .A(Red_AddKeyXOR1_XORInst_2_0_n1), 
        .B(Red_SelectedKey[42]), .ZN(Red_final[42]) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_2_0_U1 ( .A(1'b0), .B(Red_MCOutput[42]), 
        .ZN(Red_AddKeyXOR1_XORInst_2_0_n1) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_2_1_U2 ( .A(Red_AddKeyXOR1_XORInst_2_1_n1), 
        .B(Red_SelectedKey[43]), .ZN(Red_final[43]) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_2_1_U1 ( .A(1'b0), .B(Red_MCOutput[43]), 
        .ZN(Red_AddKeyXOR1_XORInst_2_1_n1) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_2_2_U2 ( .A(Red_AddKeyXOR1_XORInst_2_2_n1), 
        .B(Red_SelectedKey[44]), .ZN(Red_final[44]) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_2_2_U1 ( .A(1'b0), .B(Red_MCOutput[44]), 
        .ZN(Red_AddKeyXOR1_XORInst_2_2_n1) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_3_0_U2 ( .A(Red_AddKeyXOR1_XORInst_3_0_n1), 
        .B(Red_SelectedKey[45]), .ZN(Red_final[45]) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_3_0_U1 ( .A(1'b0), .B(Red_MCOutput[45]), 
        .ZN(Red_AddKeyXOR1_XORInst_3_0_n1) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_3_1_U2 ( .A(Red_AddKeyXOR1_XORInst_3_1_n1), 
        .B(Red_SelectedKey[46]), .ZN(Red_final[46]) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_3_1_U1 ( .A(1'b0), .B(Red_MCOutput[46]), 
        .ZN(Red_AddKeyXOR1_XORInst_3_1_n1) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_3_2_U2 ( .A(Red_AddKeyXOR1_XORInst_3_2_n1), 
        .B(Red_SelectedKey[47]), .ZN(Red_final[47]) );
  XNOR2_X1 Red_AddKeyXOR1_XORInst_3_2_U1 ( .A(1'b0), .B(Red_MCOutput[47]), 
        .ZN(Red_AddKeyXOR1_XORInst_3_2_n1) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_0_U3 ( .A(
        Red_AddKeyConstXOR_XORInst_0_0_n2), .B(
        Red_AddKeyConstXOR_XORInst_0_0_n1), .ZN(Red_final[30]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_0_U2 ( .A(Red_SelectedKey[30]), .B(
        Red_RoundConstant[0]), .ZN(Red_AddKeyConstXOR_XORInst_0_0_n1) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_0_0_U1 ( .A(1'b0), .B(Red_MCOutput[30]), 
        .Z(Red_AddKeyConstXOR_XORInst_0_0_n2) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_1_U3 ( .A(
        Red_AddKeyConstXOR_XORInst_0_1_n2), .B(
        Red_AddKeyConstXOR_XORInst_0_1_n1), .ZN(Red_final[31]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_1_U2 ( .A(Red_SelectedKey[31]), .B(
        Red_RoundConstant[1]), .ZN(Red_AddKeyConstXOR_XORInst_0_1_n1) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_0_1_U1 ( .A(1'b0), .B(Red_MCOutput[31]), 
        .Z(Red_AddKeyConstXOR_XORInst_0_1_n2) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_2_U3 ( .A(
        Red_AddKeyConstXOR_XORInst_0_2_n2), .B(
        Red_AddKeyConstXOR_XORInst_0_2_n1), .ZN(Red_final[32]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_0_2_U2 ( .A(Red_SelectedKey[32]), .B(
        Red_RoundConstant[2]), .ZN(Red_AddKeyConstXOR_XORInst_0_2_n1) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_0_2_U1 ( .A(1'b0), .B(Red_MCOutput[32]), 
        .Z(Red_AddKeyConstXOR_XORInst_0_2_n2) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_0_U3 ( .A(
        Red_AddKeyConstXOR_XORInst_1_0_n2), .B(
        Red_AddKeyConstXOR_XORInst_1_0_n1), .ZN(Red_final[33]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_0_U2 ( .A(Red_SelectedKey[33]), .B(
        Red_RoundConstant[3]), .ZN(Red_AddKeyConstXOR_XORInst_1_0_n1) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_1_0_U1 ( .A(1'b0), .B(Red_MCOutput[33]), 
        .Z(Red_AddKeyConstXOR_XORInst_1_0_n2) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_1_U3 ( .A(
        Red_AddKeyConstXOR_XORInst_1_1_n2), .B(
        Red_AddKeyConstXOR_XORInst_1_1_n1), .ZN(Red_final[34]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_1_U2 ( .A(Red_SelectedKey[34]), .B(
        Red_RoundConstant[4]), .ZN(Red_AddKeyConstXOR_XORInst_1_1_n1) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_1_1_U1 ( .A(1'b0), .B(Red_MCOutput[34]), 
        .Z(Red_AddKeyConstXOR_XORInst_1_1_n2) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_2_U3 ( .A(
        Red_AddKeyConstXOR_XORInst_1_2_n2), .B(
        Red_AddKeyConstXOR_XORInst_1_2_n1), .ZN(Red_final[35]) );
  XNOR2_X1 Red_AddKeyConstXOR_XORInst_1_2_U2 ( .A(Red_SelectedKey[35]), .B(
        Red_RoundConstant[5]), .ZN(Red_AddKeyConstXOR_XORInst_1_2_n1) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_1_2_U1 ( .A(1'b0), .B(Red_MCOutput[35]), 
        .Z(Red_AddKeyConstXOR_XORInst_1_2_n2) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_0_0_U2 ( .A(Red_AddKeyXOR2_XORInst_0_0_n1), 
        .B(Red_SelectedKey[0]), .ZN(Red_final[0]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_0_0_U1 ( .A(1'b0), .B(Red_MCOutput[0]), .ZN(
        Red_AddKeyXOR2_XORInst_0_0_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_0_1_U2 ( .A(Red_AddKeyXOR2_XORInst_0_1_n1), 
        .B(Red_SelectedKey[1]), .ZN(Red_final[1]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_0_1_U1 ( .A(1'b0), .B(Red_MCOutput[1]), .ZN(
        Red_AddKeyXOR2_XORInst_0_1_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_0_2_U2 ( .A(Red_AddKeyXOR2_XORInst_0_2_n1), 
        .B(Red_SelectedKey[2]), .ZN(Red_final[2]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_0_2_U1 ( .A(1'b0), .B(Red_MCOutput[2]), .ZN(
        Red_AddKeyXOR2_XORInst_0_2_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_1_0_U2 ( .A(Red_AddKeyXOR2_XORInst_1_0_n1), 
        .B(Red_SelectedKey[3]), .ZN(Red_final[3]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_1_0_U1 ( .A(1'b0), .B(Red_MCOutput[3]), .ZN(
        Red_AddKeyXOR2_XORInst_1_0_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_1_1_U2 ( .A(Red_AddKeyXOR2_XORInst_1_1_n1), 
        .B(Red_SelectedKey[4]), .ZN(Red_final[4]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_1_1_U1 ( .A(1'b0), .B(Red_MCOutput[4]), .ZN(
        Red_AddKeyXOR2_XORInst_1_1_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_1_2_U2 ( .A(Red_AddKeyXOR2_XORInst_1_2_n1), 
        .B(Red_SelectedKey[5]), .ZN(Red_final[5]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_1_2_U1 ( .A(1'b0), .B(Red_MCOutput[5]), .ZN(
        Red_AddKeyXOR2_XORInst_1_2_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_2_0_U2 ( .A(Red_AddKeyXOR2_XORInst_2_0_n1), 
        .B(Red_SelectedKey[6]), .ZN(Red_final[6]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_2_0_U1 ( .A(1'b0), .B(Red_MCOutput[6]), .ZN(
        Red_AddKeyXOR2_XORInst_2_0_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_2_1_U2 ( .A(Red_AddKeyXOR2_XORInst_2_1_n1), 
        .B(Red_SelectedKey[7]), .ZN(Red_final[7]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_2_1_U1 ( .A(1'b0), .B(Red_MCOutput[7]), .ZN(
        Red_AddKeyXOR2_XORInst_2_1_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_2_2_U2 ( .A(Red_AddKeyXOR2_XORInst_2_2_n1), 
        .B(Red_SelectedKey[8]), .ZN(Red_final[8]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_2_2_U1 ( .A(1'b0), .B(Red_MCOutput[8]), .ZN(
        Red_AddKeyXOR2_XORInst_2_2_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_3_0_U2 ( .A(Red_AddKeyXOR2_XORInst_3_0_n1), 
        .B(Red_SelectedKey[9]), .ZN(Red_final[9]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_3_0_U1 ( .A(1'b0), .B(Red_MCOutput[9]), .ZN(
        Red_AddKeyXOR2_XORInst_3_0_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_3_1_U2 ( .A(Red_AddKeyXOR2_XORInst_3_1_n1), 
        .B(Red_SelectedKey[10]), .ZN(Red_final[10]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_3_1_U1 ( .A(1'b0), .B(Red_MCOutput[10]), 
        .ZN(Red_AddKeyXOR2_XORInst_3_1_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_3_2_U2 ( .A(Red_AddKeyXOR2_XORInst_3_2_n1), 
        .B(Red_SelectedKey[11]), .ZN(Red_final[11]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_3_2_U1 ( .A(1'b0), .B(Red_MCOutput[11]), 
        .ZN(Red_AddKeyXOR2_XORInst_3_2_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_4_0_U2 ( .A(Red_AddKeyXOR2_XORInst_4_0_n1), 
        .B(Red_SelectedKey[12]), .ZN(Red_final[12]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_4_0_U1 ( .A(1'b0), .B(Red_MCOutput[12]), 
        .ZN(Red_AddKeyXOR2_XORInst_4_0_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_4_1_U2 ( .A(Red_AddKeyXOR2_XORInst_4_1_n1), 
        .B(Red_SelectedKey[13]), .ZN(Red_final[13]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_4_1_U1 ( .A(1'b0), .B(Red_MCOutput[13]), 
        .ZN(Red_AddKeyXOR2_XORInst_4_1_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_4_2_U2 ( .A(Red_AddKeyXOR2_XORInst_4_2_n1), 
        .B(Red_SelectedKey[14]), .ZN(Red_final[14]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_4_2_U1 ( .A(1'b0), .B(Red_MCOutput[14]), 
        .ZN(Red_AddKeyXOR2_XORInst_4_2_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_5_0_U2 ( .A(Red_AddKeyXOR2_XORInst_5_0_n1), 
        .B(Red_SelectedKey[15]), .ZN(Red_final[15]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_5_0_U1 ( .A(1'b0), .B(Red_MCOutput[15]), 
        .ZN(Red_AddKeyXOR2_XORInst_5_0_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_5_1_U2 ( .A(Red_AddKeyXOR2_XORInst_5_1_n1), 
        .B(Red_SelectedKey[16]), .ZN(Red_final[16]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_5_1_U1 ( .A(1'b0), .B(Red_MCOutput[16]), 
        .ZN(Red_AddKeyXOR2_XORInst_5_1_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_5_2_U2 ( .A(Red_AddKeyXOR2_XORInst_5_2_n1), 
        .B(Red_SelectedKey[17]), .ZN(Red_final[17]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_5_2_U1 ( .A(1'b0), .B(Red_MCOutput[17]), 
        .ZN(Red_AddKeyXOR2_XORInst_5_2_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_6_0_U2 ( .A(Red_AddKeyXOR2_XORInst_6_0_n1), 
        .B(Red_SelectedKey[18]), .ZN(Red_final[18]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_6_0_U1 ( .A(1'b0), .B(Red_MCOutput[18]), 
        .ZN(Red_AddKeyXOR2_XORInst_6_0_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_6_1_U2 ( .A(Red_AddKeyXOR2_XORInst_6_1_n1), 
        .B(Red_SelectedKey[19]), .ZN(Red_final[19]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_6_1_U1 ( .A(1'b0), .B(Red_MCOutput[19]), 
        .ZN(Red_AddKeyXOR2_XORInst_6_1_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_6_2_U2 ( .A(Red_AddKeyXOR2_XORInst_6_2_n1), 
        .B(Red_SelectedKey[20]), .ZN(Red_final[20]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_6_2_U1 ( .A(1'b0), .B(Red_MCOutput[20]), 
        .ZN(Red_AddKeyXOR2_XORInst_6_2_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_7_0_U2 ( .A(Red_AddKeyXOR2_XORInst_7_0_n1), 
        .B(Red_SelectedKey[21]), .ZN(Red_final[21]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_7_0_U1 ( .A(1'b0), .B(Red_MCOutput[21]), 
        .ZN(Red_AddKeyXOR2_XORInst_7_0_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_7_1_U2 ( .A(Red_AddKeyXOR2_XORInst_7_1_n1), 
        .B(Red_SelectedKey[22]), .ZN(Red_final[22]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_7_1_U1 ( .A(1'b0), .B(Red_MCOutput[22]), 
        .ZN(Red_AddKeyXOR2_XORInst_7_1_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_7_2_U2 ( .A(Red_AddKeyXOR2_XORInst_7_2_n1), 
        .B(Red_SelectedKey[23]), .ZN(Red_final[23]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_7_2_U1 ( .A(1'b0), .B(Red_MCOutput[23]), 
        .ZN(Red_AddKeyXOR2_XORInst_7_2_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_8_0_U2 ( .A(Red_AddKeyXOR2_XORInst_8_0_n1), 
        .B(Red_SelectedKey[24]), .ZN(Red_final[24]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_8_0_U1 ( .A(1'b0), .B(Red_MCOutput[24]), 
        .ZN(Red_AddKeyXOR2_XORInst_8_0_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_8_1_U2 ( .A(Red_AddKeyXOR2_XORInst_8_1_n1), 
        .B(Red_SelectedKey[25]), .ZN(Red_final[25]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_8_1_U1 ( .A(1'b0), .B(Red_MCOutput[25]), 
        .ZN(Red_AddKeyXOR2_XORInst_8_1_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_8_2_U2 ( .A(Red_AddKeyXOR2_XORInst_8_2_n1), 
        .B(Red_SelectedKey[26]), .ZN(Red_final[26]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_8_2_U1 ( .A(1'b0), .B(Red_MCOutput[26]), 
        .ZN(Red_AddKeyXOR2_XORInst_8_2_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_9_0_U2 ( .A(Red_AddKeyXOR2_XORInst_9_0_n1), 
        .B(Red_SelectedKey[27]), .ZN(Red_final[27]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_9_0_U1 ( .A(1'b0), .B(Red_MCOutput[27]), 
        .ZN(Red_AddKeyXOR2_XORInst_9_0_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_9_1_U2 ( .A(Red_AddKeyXOR2_XORInst_9_1_n1), 
        .B(Red_SelectedKey[28]), .ZN(Red_final[28]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_9_1_U1 ( .A(1'b0), .B(Red_MCOutput[28]), 
        .ZN(Red_AddKeyXOR2_XORInst_9_1_n1) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_9_2_U2 ( .A(Red_AddKeyXOR2_XORInst_9_2_n1), 
        .B(Red_SelectedKey[29]), .ZN(Red_final[29]) );
  XNOR2_X1 Red_AddKeyXOR2_XORInst_9_2_U1 ( .A(1'b0), .B(Red_MCOutput[29]), 
        .ZN(Red_AddKeyXOR2_XORInst_9_2_n1) );
  DFF_X1 Red_StateReg_s_current_state_reg_0_ ( .D(Red_final[0]), .CK(clk), .Q(
        Red_StateRegOutput[0]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_1_ ( .D(Red_final[1]), .CK(clk), .Q(
        Red_StateRegOutput[1]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_2_ ( .D(Red_final[2]), .CK(clk), .Q(
        Red_StateRegOutput[2]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_3_ ( .D(Red_final[3]), .CK(clk), .Q(
        Red_StateRegOutput[3]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_4_ ( .D(Red_final[4]), .CK(clk), .Q(
        Red_StateRegOutput[4]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_5_ ( .D(Red_final[5]), .CK(clk), .Q(
        Red_StateRegOutput[5]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_6_ ( .D(Red_final[6]), .CK(clk), .Q(
        Red_StateRegOutput[6]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_7_ ( .D(Red_final[7]), .CK(clk), .Q(
        Red_StateRegOutput[7]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_8_ ( .D(Red_final[8]), .CK(clk), .Q(
        Red_StateRegOutput[8]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_9_ ( .D(Red_final[9]), .CK(clk), .Q(
        Red_StateRegOutput[9]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_10_ ( .D(Red_final[10]), .CK(clk), 
        .Q(Red_StateRegOutput[10]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_11_ ( .D(Red_final[11]), .CK(clk), 
        .Q(Red_StateRegOutput[11]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_12_ ( .D(Red_final[12]), .CK(clk), 
        .Q(Red_StateRegOutput[12]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_13_ ( .D(Red_final[13]), .CK(clk), 
        .Q(Red_StateRegOutput[13]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_14_ ( .D(Red_final[14]), .CK(clk), 
        .Q(Red_StateRegOutput[14]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_15_ ( .D(Red_final[15]), .CK(clk), 
        .Q(Red_StateRegOutput[15]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_16_ ( .D(Red_final[16]), .CK(clk), 
        .Q(Red_StateRegOutput[16]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_17_ ( .D(Red_final[17]), .CK(clk), 
        .Q(Red_StateRegOutput[17]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_18_ ( .D(Red_final[18]), .CK(clk), 
        .Q(Red_StateRegOutput[18]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_19_ ( .D(Red_final[19]), .CK(clk), 
        .Q(Red_StateRegOutput[19]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_20_ ( .D(Red_final[20]), .CK(clk), 
        .Q(Red_StateRegOutput[20]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_21_ ( .D(Red_final[21]), .CK(clk), 
        .Q(Red_StateRegOutput[21]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_22_ ( .D(Red_final[22]), .CK(clk), 
        .Q(Red_StateRegOutput[22]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_23_ ( .D(Red_final[23]), .CK(clk), 
        .Q(Red_StateRegOutput[23]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_24_ ( .D(Red_final[24]), .CK(clk), 
        .Q(Red_StateRegOutput[24]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_25_ ( .D(Red_final[25]), .CK(clk), 
        .Q(Red_StateRegOutput[25]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_26_ ( .D(Red_final[26]), .CK(clk), 
        .Q(Red_StateRegOutput[26]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_27_ ( .D(Red_final[27]), .CK(clk), 
        .Q(Red_StateRegOutput[27]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_28_ ( .D(Red_final[28]), .CK(clk), 
        .Q(Red_StateRegOutput[28]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_29_ ( .D(Red_final[29]), .CK(clk), 
        .Q(Red_StateRegOutput[29]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_30_ ( .D(Red_final[30]), .CK(clk), 
        .Q(Red_StateRegOutput[30]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_31_ ( .D(Red_final[31]), .CK(clk), 
        .Q(Red_StateRegOutput[31]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_32_ ( .D(Red_final[32]), .CK(clk), 
        .Q(Red_StateRegOutput[32]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_33_ ( .D(Red_final[33]), .CK(clk), 
        .Q(Red_StateRegOutput[33]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_34_ ( .D(Red_final[34]), .CK(clk), 
        .Q(Red_StateRegOutput[34]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_35_ ( .D(Red_final[35]), .CK(clk), 
        .Q(Red_StateRegOutput[35]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_36_ ( .D(Red_final[36]), .CK(clk), 
        .Q(Red_StateRegOutput[36]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_37_ ( .D(Red_final[37]), .CK(clk), 
        .Q(Red_StateRegOutput[37]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_38_ ( .D(Red_final[38]), .CK(clk), 
        .Q(Red_StateRegOutput[38]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_39_ ( .D(Red_final[39]), .CK(clk), 
        .Q(Red_StateRegOutput[39]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_40_ ( .D(Red_final[40]), .CK(clk), 
        .Q(Red_StateRegOutput[40]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_41_ ( .D(Red_final[41]), .CK(clk), 
        .Q(Red_StateRegOutput[41]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_42_ ( .D(Red_final[42]), .CK(clk), 
        .Q(Red_StateRegOutput[42]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_43_ ( .D(Red_final[43]), .CK(clk), 
        .Q(Red_StateRegOutput[43]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_44_ ( .D(Red_final[44]), .CK(clk), 
        .Q(Red_StateRegOutput[44]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_45_ ( .D(Red_final[45]), .CK(clk), 
        .Q(Red_StateRegOutput[45]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_46_ ( .D(Red_final[46]), .CK(clk), 
        .Q(Red_StateRegOutput[46]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_47_ ( .D(Red_final[47]), .CK(clk), 
        .Q(Red_StateRegOutput[47]), .QN() );
  XOR2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U3 ( .A(PermutationOutput[1]), .B(
        Red_SubCellInst_LFInst_0_LFInst_0_n2), .Z(Red_Feedback[0]) );
  OAI21_X1 Red_SubCellInst_LFInst_0_LFInst_0_U2 ( .B1(PermutationOutput[3]), 
        .B2(PermutationOutput[2]), .A(Red_SubCellInst_LFInst_0_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_0_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U1 ( .A1(PermutationOutput[3]), 
        .A2(PermutationOutput[0]), .ZN(Red_SubCellInst_LFInst_0_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_0_LFInst_1_U5 ( .A1(PermutationOutput[0]), 
        .A2(Red_SubCellInst_LFInst_0_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_0_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_0_LFInst_1_n2), .ZN(Red_Feedback[1]) );
  OAI21_X1 Red_SubCellInst_LFInst_0_LFInst_1_U4 ( .B1(PermutationOutput[1]), 
        .B2(PermutationOutput[2]), .A(PermutationOutput[0]), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_0_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_0_LFInst_1_n2), .B(PermutationOutput[2]), .Z(
        Red_SubCellInst_LFInst_0_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_0_LFInst_1_U2 ( .A1(PermutationOutput[3]), 
        .A2(Red_SubCellInst_LFInst_0_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_0_LFInst_1_U1 ( .A(PermutationOutput[1]), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_0_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_0_LFInst_2_n6), .B2(PermutationOutput[2]), .C1(
        Red_SubCellInst_LFInst_0_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_0_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_0_LFInst_2_n3), .ZN(Red_Feedback[2]) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_0_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U5 ( .A1(PermutationOutput[1]), 
        .A2(Red_SubCellInst_LFInst_0_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_0_LFInst_2_U4 ( .A(PermutationOutput[3]), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U3 ( .A1(PermutationOutput[2]), 
        .A2(Red_SubCellInst_LFInst_0_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_0_LFInst_2_U2 ( .A(PermutationOutput[0]), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_2_U1 ( .A1(PermutationOutput[1]), 
        .A2(PermutationOutput[0]), .ZN(Red_SubCellInst_LFInst_0_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U3 ( .A(PermutationOutput[5]), .B(
        Red_SubCellInst_LFInst_1_LFInst_0_n2), .Z(Red_Feedback[3]) );
  OAI21_X1 Red_SubCellInst_LFInst_1_LFInst_0_U2 ( .B1(PermutationOutput[7]), 
        .B2(PermutationOutput[6]), .A(Red_SubCellInst_LFInst_1_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_1_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U1 ( .A1(PermutationOutput[7]), 
        .A2(PermutationOutput[4]), .ZN(Red_SubCellInst_LFInst_1_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_1_LFInst_1_U5 ( .A1(PermutationOutput[4]), 
        .A2(Red_SubCellInst_LFInst_1_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_1_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_1_LFInst_1_n2), .ZN(Red_Feedback[4]) );
  OAI21_X1 Red_SubCellInst_LFInst_1_LFInst_1_U4 ( .B1(PermutationOutput[5]), 
        .B2(PermutationOutput[6]), .A(PermutationOutput[4]), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_1_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_1_LFInst_1_n2), .B(PermutationOutput[6]), .Z(
        Red_SubCellInst_LFInst_1_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_1_LFInst_1_U2 ( .A1(PermutationOutput[7]), 
        .A2(Red_SubCellInst_LFInst_1_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_1_LFInst_1_U1 ( .A(PermutationOutput[5]), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_1_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_1_LFInst_2_n6), .B2(PermutationOutput[6]), .C1(
        Red_SubCellInst_LFInst_1_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_1_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_1_LFInst_2_n3), .ZN(Red_Feedback[5]) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_1_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U5 ( .A1(PermutationOutput[5]), 
        .A2(Red_SubCellInst_LFInst_1_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_1_LFInst_2_U4 ( .A(PermutationOutput[7]), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U3 ( .A1(PermutationOutput[6]), 
        .A2(Red_SubCellInst_LFInst_1_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_1_LFInst_2_U2 ( .A(PermutationOutput[4]), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_2_U1 ( .A1(PermutationOutput[5]), 
        .A2(PermutationOutput[4]), .ZN(Red_SubCellInst_LFInst_1_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U3 ( .A(PermutationOutput[9]), .B(
        Red_SubCellInst_LFInst_2_LFInst_0_n2), .Z(Red_Feedback[6]) );
  OAI21_X1 Red_SubCellInst_LFInst_2_LFInst_0_U2 ( .B1(PermutationOutput[11]), 
        .B2(PermutationOutput[10]), .A(Red_SubCellInst_LFInst_2_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U1 ( .A1(PermutationOutput[11]), 
        .A2(PermutationOutput[8]), .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_2_LFInst_1_U5 ( .A1(PermutationOutput[8]), 
        .A2(Red_SubCellInst_LFInst_2_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_2_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_2_LFInst_1_n2), .ZN(Red_Feedback[7]) );
  OAI21_X1 Red_SubCellInst_LFInst_2_LFInst_1_U4 ( .B1(PermutationOutput[9]), 
        .B2(PermutationOutput[10]), .A(PermutationOutput[8]), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_2_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_2_LFInst_1_n2), .B(PermutationOutput[10]), .Z(
        Red_SubCellInst_LFInst_2_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_2_LFInst_1_U2 ( .A1(PermutationOutput[11]), 
        .A2(Red_SubCellInst_LFInst_2_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_2_LFInst_1_U1 ( .A(PermutationOutput[9]), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_2_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_2_LFInst_2_n6), .B2(PermutationOutput[10]), 
        .C1(Red_SubCellInst_LFInst_2_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_2_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_2_LFInst_2_n3), .ZN(Red_Feedback[8]) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_2_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U5 ( .A1(PermutationOutput[9]), 
        .A2(Red_SubCellInst_LFInst_2_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_2_LFInst_2_U4 ( .A(PermutationOutput[11]), 
        .ZN(Red_SubCellInst_LFInst_2_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U3 ( .A1(PermutationOutput[10]), 
        .A2(Red_SubCellInst_LFInst_2_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_2_LFInst_2_U2 ( .A(PermutationOutput[8]), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_2_U1 ( .A1(PermutationOutput[9]), 
        .A2(PermutationOutput[8]), .ZN(Red_SubCellInst_LFInst_2_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U3 ( .A(PermutationOutput[13]), 
        .B(Red_SubCellInst_LFInst_3_LFInst_0_n2), .Z(Red_Feedback[9]) );
  OAI21_X1 Red_SubCellInst_LFInst_3_LFInst_0_U2 ( .B1(PermutationOutput[15]), 
        .B2(PermutationOutput[14]), .A(Red_SubCellInst_LFInst_3_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U1 ( .A1(PermutationOutput[15]), 
        .A2(PermutationOutput[12]), .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_3_LFInst_1_U5 ( .A1(PermutationOutput[12]), 
        .A2(Red_SubCellInst_LFInst_3_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_3_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_3_LFInst_1_n2), .ZN(Red_Feedback[10]) );
  OAI21_X1 Red_SubCellInst_LFInst_3_LFInst_1_U4 ( .B1(PermutationOutput[13]), 
        .B2(PermutationOutput[14]), .A(PermutationOutput[12]), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_3_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_3_LFInst_1_n2), .B(PermutationOutput[14]), .Z(
        Red_SubCellInst_LFInst_3_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_3_LFInst_1_U2 ( .A1(PermutationOutput[15]), 
        .A2(Red_SubCellInst_LFInst_3_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_3_LFInst_1_U1 ( .A(PermutationOutput[13]), 
        .ZN(Red_SubCellInst_LFInst_3_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_3_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_3_LFInst_2_n6), .B2(PermutationOutput[14]), 
        .C1(Red_SubCellInst_LFInst_3_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_3_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_3_LFInst_2_n3), .ZN(Red_Feedback[11]) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_3_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U5 ( .A1(PermutationOutput[13]), 
        .A2(Red_SubCellInst_LFInst_3_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_3_LFInst_2_U4 ( .A(PermutationOutput[15]), 
        .ZN(Red_SubCellInst_LFInst_3_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U3 ( .A1(PermutationOutput[14]), 
        .A2(Red_SubCellInst_LFInst_3_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_3_LFInst_2_U2 ( .A(PermutationOutput[12]), 
        .ZN(Red_SubCellInst_LFInst_3_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_2_U1 ( .A1(PermutationOutput[13]), 
        .A2(PermutationOutput[12]), .ZN(Red_SubCellInst_LFInst_3_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U3 ( .A(PermutationOutput[17]), 
        .B(Red_SubCellInst_LFInst_4_LFInst_0_n2), .Z(Red_Feedback[12]) );
  OAI21_X1 Red_SubCellInst_LFInst_4_LFInst_0_U2 ( .B1(PermutationOutput[19]), 
        .B2(PermutationOutput[18]), .A(Red_SubCellInst_LFInst_4_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U1 ( .A1(PermutationOutput[19]), 
        .A2(PermutationOutput[16]), .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_4_LFInst_1_U5 ( .A1(PermutationOutput[16]), 
        .A2(Red_SubCellInst_LFInst_4_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_4_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_4_LFInst_1_n2), .ZN(Red_Feedback[13]) );
  OAI21_X1 Red_SubCellInst_LFInst_4_LFInst_1_U4 ( .B1(PermutationOutput[17]), 
        .B2(PermutationOutput[18]), .A(PermutationOutput[16]), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_4_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_4_LFInst_1_n2), .B(PermutationOutput[18]), .Z(
        Red_SubCellInst_LFInst_4_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_4_LFInst_1_U2 ( .A1(PermutationOutput[19]), 
        .A2(Red_SubCellInst_LFInst_4_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_4_LFInst_1_U1 ( .A(PermutationOutput[17]), 
        .ZN(Red_SubCellInst_LFInst_4_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_4_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_4_LFInst_2_n6), .B2(PermutationOutput[18]), 
        .C1(Red_SubCellInst_LFInst_4_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_4_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_4_LFInst_2_n3), .ZN(Red_Feedback[14]) );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_4_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U5 ( .A1(PermutationOutput[17]), 
        .A2(Red_SubCellInst_LFInst_4_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_4_LFInst_2_U4 ( .A(PermutationOutput[19]), 
        .ZN(Red_SubCellInst_LFInst_4_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U3 ( .A1(PermutationOutput[18]), 
        .A2(Red_SubCellInst_LFInst_4_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_4_LFInst_2_U2 ( .A(PermutationOutput[16]), 
        .ZN(Red_SubCellInst_LFInst_4_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_2_U1 ( .A1(PermutationOutput[17]), 
        .A2(PermutationOutput[16]), .ZN(Red_SubCellInst_LFInst_4_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U3 ( .A(PermutationOutput[21]), 
        .B(Red_SubCellInst_LFInst_5_LFInst_0_n2), .Z(Red_Feedback[15]) );
  OAI21_X1 Red_SubCellInst_LFInst_5_LFInst_0_U2 ( .B1(PermutationOutput[23]), 
        .B2(PermutationOutput[22]), .A(Red_SubCellInst_LFInst_5_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U1 ( .A1(PermutationOutput[23]), 
        .A2(PermutationOutput[20]), .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_5_LFInst_1_U5 ( .A1(PermutationOutput[20]), 
        .A2(Red_SubCellInst_LFInst_5_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_5_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_5_LFInst_1_n2), .ZN(Red_Feedback[16]) );
  OAI21_X1 Red_SubCellInst_LFInst_5_LFInst_1_U4 ( .B1(PermutationOutput[21]), 
        .B2(PermutationOutput[22]), .A(PermutationOutput[20]), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_5_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_5_LFInst_1_n2), .B(PermutationOutput[22]), .Z(
        Red_SubCellInst_LFInst_5_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_5_LFInst_1_U2 ( .A1(PermutationOutput[23]), 
        .A2(Red_SubCellInst_LFInst_5_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_5_LFInst_1_U1 ( .A(PermutationOutput[21]), 
        .ZN(Red_SubCellInst_LFInst_5_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_5_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_5_LFInst_2_n6), .B2(PermutationOutput[22]), 
        .C1(Red_SubCellInst_LFInst_5_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_5_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_5_LFInst_2_n3), .ZN(Red_Feedback[17]) );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_5_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U5 ( .A1(PermutationOutput[21]), 
        .A2(Red_SubCellInst_LFInst_5_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_5_LFInst_2_U4 ( .A(PermutationOutput[23]), 
        .ZN(Red_SubCellInst_LFInst_5_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U3 ( .A1(PermutationOutput[22]), 
        .A2(Red_SubCellInst_LFInst_5_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_5_LFInst_2_U2 ( .A(PermutationOutput[20]), 
        .ZN(Red_SubCellInst_LFInst_5_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_2_U1 ( .A1(PermutationOutput[21]), 
        .A2(PermutationOutput[20]), .ZN(Red_SubCellInst_LFInst_5_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U3 ( .A(PermutationOutput[25]), 
        .B(Red_SubCellInst_LFInst_6_LFInst_0_n2), .Z(Red_Feedback[18]) );
  OAI21_X1 Red_SubCellInst_LFInst_6_LFInst_0_U2 ( .B1(PermutationOutput[27]), 
        .B2(PermutationOutput[26]), .A(Red_SubCellInst_LFInst_6_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U1 ( .A1(PermutationOutput[27]), 
        .A2(PermutationOutput[24]), .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_6_LFInst_1_U5 ( .A1(PermutationOutput[24]), 
        .A2(Red_SubCellInst_LFInst_6_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_6_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_6_LFInst_1_n2), .ZN(Red_Feedback[19]) );
  OAI21_X1 Red_SubCellInst_LFInst_6_LFInst_1_U4 ( .B1(PermutationOutput[25]), 
        .B2(PermutationOutput[26]), .A(PermutationOutput[24]), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_6_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_6_LFInst_1_n2), .B(PermutationOutput[26]), .Z(
        Red_SubCellInst_LFInst_6_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_6_LFInst_1_U2 ( .A1(PermutationOutput[27]), 
        .A2(Red_SubCellInst_LFInst_6_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_6_LFInst_1_U1 ( .A(PermutationOutput[25]), 
        .ZN(Red_SubCellInst_LFInst_6_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_6_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_6_LFInst_2_n6), .B2(PermutationOutput[26]), 
        .C1(Red_SubCellInst_LFInst_6_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_6_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_6_LFInst_2_n3), .ZN(Red_Feedback[20]) );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_6_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U5 ( .A1(PermutationOutput[25]), 
        .A2(Red_SubCellInst_LFInst_6_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_6_LFInst_2_U4 ( .A(PermutationOutput[27]), 
        .ZN(Red_SubCellInst_LFInst_6_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U3 ( .A1(PermutationOutput[26]), 
        .A2(Red_SubCellInst_LFInst_6_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_6_LFInst_2_U2 ( .A(PermutationOutput[24]), 
        .ZN(Red_SubCellInst_LFInst_6_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_2_U1 ( .A1(PermutationOutput[25]), 
        .A2(PermutationOutput[24]), .ZN(Red_SubCellInst_LFInst_6_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U3 ( .A(PermutationOutput[29]), 
        .B(Red_SubCellInst_LFInst_7_LFInst_0_n2), .Z(Red_Feedback[21]) );
  OAI21_X1 Red_SubCellInst_LFInst_7_LFInst_0_U2 ( .B1(PermutationOutput[31]), 
        .B2(PermutationOutput[30]), .A(Red_SubCellInst_LFInst_7_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U1 ( .A1(PermutationOutput[31]), 
        .A2(PermutationOutput[28]), .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_7_LFInst_1_U5 ( .A1(PermutationOutput[28]), 
        .A2(Red_SubCellInst_LFInst_7_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_7_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_7_LFInst_1_n2), .ZN(Red_Feedback[22]) );
  OAI21_X1 Red_SubCellInst_LFInst_7_LFInst_1_U4 ( .B1(PermutationOutput[29]), 
        .B2(PermutationOutput[30]), .A(PermutationOutput[28]), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_7_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_7_LFInst_1_n2), .B(PermutationOutput[30]), .Z(
        Red_SubCellInst_LFInst_7_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_7_LFInst_1_U2 ( .A1(PermutationOutput[31]), 
        .A2(Red_SubCellInst_LFInst_7_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_7_LFInst_1_U1 ( .A(PermutationOutput[29]), 
        .ZN(Red_SubCellInst_LFInst_7_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_7_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_7_LFInst_2_n6), .B2(PermutationOutput[30]), 
        .C1(Red_SubCellInst_LFInst_7_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_7_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_7_LFInst_2_n3), .ZN(Red_Feedback[23]) );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_7_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U5 ( .A1(PermutationOutput[29]), 
        .A2(Red_SubCellInst_LFInst_7_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_7_LFInst_2_U4 ( .A(PermutationOutput[31]), 
        .ZN(Red_SubCellInst_LFInst_7_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U3 ( .A1(PermutationOutput[30]), 
        .A2(Red_SubCellInst_LFInst_7_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_7_LFInst_2_U2 ( .A(PermutationOutput[28]), 
        .ZN(Red_SubCellInst_LFInst_7_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_2_U1 ( .A1(PermutationOutput[29]), 
        .A2(PermutationOutput[28]), .ZN(Red_SubCellInst_LFInst_7_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U3 ( .A(PermutationOutput[33]), 
        .B(Red_SubCellInst_LFInst_8_LFInst_0_n2), .Z(Red_Feedback[24]) );
  OAI21_X1 Red_SubCellInst_LFInst_8_LFInst_0_U2 ( .B1(PermutationOutput[35]), 
        .B2(PermutationOutput[34]), .A(Red_SubCellInst_LFInst_8_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U1 ( .A1(PermutationOutput[35]), 
        .A2(PermutationOutput[32]), .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_8_LFInst_1_U5 ( .A1(PermutationOutput[32]), 
        .A2(Red_SubCellInst_LFInst_8_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_8_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_8_LFInst_1_n2), .ZN(Red_Feedback[25]) );
  OAI21_X1 Red_SubCellInst_LFInst_8_LFInst_1_U4 ( .B1(PermutationOutput[33]), 
        .B2(PermutationOutput[34]), .A(PermutationOutput[32]), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_8_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_8_LFInst_1_n2), .B(PermutationOutput[34]), .Z(
        Red_SubCellInst_LFInst_8_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_8_LFInst_1_U2 ( .A1(PermutationOutput[35]), 
        .A2(Red_SubCellInst_LFInst_8_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_8_LFInst_1_U1 ( .A(PermutationOutput[33]), 
        .ZN(Red_SubCellInst_LFInst_8_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_8_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_8_LFInst_2_n6), .B2(PermutationOutput[34]), 
        .C1(Red_SubCellInst_LFInst_8_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_8_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_8_LFInst_2_n3), .ZN(Red_Feedback[26]) );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_8_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U5 ( .A1(PermutationOutput[33]), 
        .A2(Red_SubCellInst_LFInst_8_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_8_LFInst_2_U4 ( .A(PermutationOutput[35]), 
        .ZN(Red_SubCellInst_LFInst_8_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U3 ( .A1(PermutationOutput[34]), 
        .A2(Red_SubCellInst_LFInst_8_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_8_LFInst_2_U2 ( .A(PermutationOutput[32]), 
        .ZN(Red_SubCellInst_LFInst_8_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_2_U1 ( .A1(PermutationOutput[33]), 
        .A2(PermutationOutput[32]), .ZN(Red_SubCellInst_LFInst_8_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U3 ( .A(PermutationOutput[37]), 
        .B(Red_SubCellInst_LFInst_9_LFInst_0_n2), .Z(Red_Feedback[27]) );
  OAI21_X1 Red_SubCellInst_LFInst_9_LFInst_0_U2 ( .B1(PermutationOutput[39]), 
        .B2(PermutationOutput[38]), .A(Red_SubCellInst_LFInst_9_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U1 ( .A1(PermutationOutput[39]), 
        .A2(PermutationOutput[36]), .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_9_LFInst_1_U5 ( .A1(PermutationOutput[36]), 
        .A2(Red_SubCellInst_LFInst_9_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_9_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_9_LFInst_1_n2), .ZN(Red_Feedback[28]) );
  OAI21_X1 Red_SubCellInst_LFInst_9_LFInst_1_U4 ( .B1(PermutationOutput[37]), 
        .B2(PermutationOutput[38]), .A(PermutationOutput[36]), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_9_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_9_LFInst_1_n2), .B(PermutationOutput[38]), .Z(
        Red_SubCellInst_LFInst_9_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_9_LFInst_1_U2 ( .A1(PermutationOutput[39]), 
        .A2(Red_SubCellInst_LFInst_9_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_9_LFInst_1_U1 ( .A(PermutationOutput[37]), 
        .ZN(Red_SubCellInst_LFInst_9_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_9_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_9_LFInst_2_n6), .B2(PermutationOutput[38]), 
        .C1(Red_SubCellInst_LFInst_9_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_9_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_9_LFInst_2_n3), .ZN(Red_Feedback[29]) );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_9_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U5 ( .A1(PermutationOutput[37]), 
        .A2(Red_SubCellInst_LFInst_9_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_9_LFInst_2_U4 ( .A(PermutationOutput[39]), 
        .ZN(Red_SubCellInst_LFInst_9_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U3 ( .A1(PermutationOutput[38]), 
        .A2(Red_SubCellInst_LFInst_9_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_9_LFInst_2_U2 ( .A(PermutationOutput[36]), 
        .ZN(Red_SubCellInst_LFInst_9_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_2_U1 ( .A1(PermutationOutput[37]), 
        .A2(PermutationOutput[36]), .ZN(Red_SubCellInst_LFInst_9_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U3 ( .A(PermutationOutput[41]), 
        .B(Red_SubCellInst_LFInst_10_LFInst_0_n2), .Z(Red_Feedback[30]) );
  OAI21_X1 Red_SubCellInst_LFInst_10_LFInst_0_U2 ( .B1(PermutationOutput[43]), 
        .B2(PermutationOutput[42]), .A(Red_SubCellInst_LFInst_10_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U1 ( .A1(PermutationOutput[43]), 
        .A2(PermutationOutput[40]), .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_10_LFInst_1_U5 ( .A1(PermutationOutput[40]), 
        .A2(Red_SubCellInst_LFInst_10_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_10_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_10_LFInst_1_n2), .ZN(Red_Feedback[31]) );
  OAI21_X1 Red_SubCellInst_LFInst_10_LFInst_1_U4 ( .B1(PermutationOutput[41]), 
        .B2(PermutationOutput[42]), .A(PermutationOutput[40]), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_10_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_10_LFInst_1_n2), .B(PermutationOutput[42]), .Z(
        Red_SubCellInst_LFInst_10_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_10_LFInst_1_U2 ( .A1(PermutationOutput[43]), 
        .A2(Red_SubCellInst_LFInst_10_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_10_LFInst_1_U1 ( .A(PermutationOutput[41]), 
        .ZN(Red_SubCellInst_LFInst_10_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_10_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_10_LFInst_2_n6), .B2(PermutationOutput[42]), 
        .C1(Red_SubCellInst_LFInst_10_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_10_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_10_LFInst_2_n3), .ZN(Red_Feedback[32]) );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_10_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U5 ( .A1(PermutationOutput[41]), 
        .A2(Red_SubCellInst_LFInst_10_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_10_LFInst_2_U4 ( .A(PermutationOutput[43]), 
        .ZN(Red_SubCellInst_LFInst_10_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U3 ( .A1(PermutationOutput[42]), 
        .A2(Red_SubCellInst_LFInst_10_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_10_LFInst_2_U2 ( .A(PermutationOutput[40]), 
        .ZN(Red_SubCellInst_LFInst_10_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_2_U1 ( .A1(PermutationOutput[41]), 
        .A2(PermutationOutput[40]), .ZN(Red_SubCellInst_LFInst_10_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U3 ( .A(PermutationOutput[45]), 
        .B(Red_SubCellInst_LFInst_11_LFInst_0_n2), .Z(Red_Feedback[33]) );
  OAI21_X1 Red_SubCellInst_LFInst_11_LFInst_0_U2 ( .B1(PermutationOutput[47]), 
        .B2(PermutationOutput[46]), .A(Red_SubCellInst_LFInst_11_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U1 ( .A1(PermutationOutput[47]), 
        .A2(PermutationOutput[44]), .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_11_LFInst_1_U5 ( .A1(PermutationOutput[44]), 
        .A2(Red_SubCellInst_LFInst_11_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_11_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_11_LFInst_1_n2), .ZN(Red_Feedback[34]) );
  OAI21_X1 Red_SubCellInst_LFInst_11_LFInst_1_U4 ( .B1(PermutationOutput[45]), 
        .B2(PermutationOutput[46]), .A(PermutationOutput[44]), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_11_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_11_LFInst_1_n2), .B(PermutationOutput[46]), .Z(
        Red_SubCellInst_LFInst_11_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_11_LFInst_1_U2 ( .A1(PermutationOutput[47]), 
        .A2(Red_SubCellInst_LFInst_11_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_11_LFInst_1_U1 ( .A(PermutationOutput[45]), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_11_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_11_LFInst_2_n6), .B2(PermutationOutput[46]), 
        .C1(Red_SubCellInst_LFInst_11_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_11_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_11_LFInst_2_n3), .ZN(Red_Feedback[35]) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_11_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U5 ( .A1(PermutationOutput[45]), 
        .A2(Red_SubCellInst_LFInst_11_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_11_LFInst_2_U4 ( .A(PermutationOutput[47]), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U3 ( .A1(PermutationOutput[46]), 
        .A2(Red_SubCellInst_LFInst_11_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_11_LFInst_2_U2 ( .A(PermutationOutput[44]), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_2_U1 ( .A1(PermutationOutput[45]), 
        .A2(PermutationOutput[44]), .ZN(Red_SubCellInst_LFInst_11_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U3 ( .A(PermutationOutput[49]), 
        .B(Red_SubCellInst_LFInst_12_LFInst_0_n2), .Z(Red_Feedback[36]) );
  OAI21_X1 Red_SubCellInst_LFInst_12_LFInst_0_U2 ( .B1(PermutationOutput[51]), 
        .B2(PermutationOutput[50]), .A(Red_SubCellInst_LFInst_12_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U1 ( .A1(PermutationOutput[51]), 
        .A2(PermutationOutput[48]), .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_12_LFInst_1_U5 ( .A1(PermutationOutput[48]), 
        .A2(Red_SubCellInst_LFInst_12_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_12_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_12_LFInst_1_n2), .ZN(Red_Feedback[37]) );
  OAI21_X1 Red_SubCellInst_LFInst_12_LFInst_1_U4 ( .B1(PermutationOutput[49]), 
        .B2(PermutationOutput[50]), .A(PermutationOutput[48]), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_12_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_12_LFInst_1_n2), .B(PermutationOutput[50]), .Z(
        Red_SubCellInst_LFInst_12_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_12_LFInst_1_U2 ( .A1(PermutationOutput[51]), 
        .A2(Red_SubCellInst_LFInst_12_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_12_LFInst_1_U1 ( .A(PermutationOutput[49]), 
        .ZN(Red_SubCellInst_LFInst_12_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_12_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_12_LFInst_2_n6), .B2(PermutationOutput[50]), 
        .C1(Red_SubCellInst_LFInst_12_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_12_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_12_LFInst_2_n3), .ZN(Red_Feedback[38]) );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_12_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U5 ( .A1(PermutationOutput[49]), 
        .A2(Red_SubCellInst_LFInst_12_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_12_LFInst_2_U4 ( .A(PermutationOutput[51]), 
        .ZN(Red_SubCellInst_LFInst_12_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U3 ( .A1(PermutationOutput[50]), 
        .A2(Red_SubCellInst_LFInst_12_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_12_LFInst_2_U2 ( .A(PermutationOutput[48]), 
        .ZN(Red_SubCellInst_LFInst_12_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_2_U1 ( .A1(PermutationOutput[49]), 
        .A2(PermutationOutput[48]), .ZN(Red_SubCellInst_LFInst_12_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U3 ( .A(PermutationOutput[53]), 
        .B(Red_SubCellInst_LFInst_13_LFInst_0_n2), .Z(Red_Feedback[39]) );
  OAI21_X1 Red_SubCellInst_LFInst_13_LFInst_0_U2 ( .B1(PermutationOutput[55]), 
        .B2(PermutationOutput[54]), .A(Red_SubCellInst_LFInst_13_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U1 ( .A1(PermutationOutput[55]), 
        .A2(PermutationOutput[52]), .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_13_LFInst_1_U5 ( .A1(PermutationOutput[52]), 
        .A2(Red_SubCellInst_LFInst_13_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_13_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_13_LFInst_1_n2), .ZN(Red_Feedback[40]) );
  OAI21_X1 Red_SubCellInst_LFInst_13_LFInst_1_U4 ( .B1(PermutationOutput[53]), 
        .B2(PermutationOutput[54]), .A(PermutationOutput[52]), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_13_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_13_LFInst_1_n2), .B(PermutationOutput[54]), .Z(
        Red_SubCellInst_LFInst_13_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_13_LFInst_1_U2 ( .A1(PermutationOutput[55]), 
        .A2(Red_SubCellInst_LFInst_13_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_13_LFInst_1_U1 ( .A(PermutationOutput[53]), 
        .ZN(Red_SubCellInst_LFInst_13_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_13_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_13_LFInst_2_n6), .B2(PermutationOutput[54]), 
        .C1(Red_SubCellInst_LFInst_13_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_13_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_13_LFInst_2_n3), .ZN(Red_Feedback[41]) );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_13_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U5 ( .A1(PermutationOutput[53]), 
        .A2(Red_SubCellInst_LFInst_13_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_13_LFInst_2_U4 ( .A(PermutationOutput[55]), 
        .ZN(Red_SubCellInst_LFInst_13_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U3 ( .A1(PermutationOutput[54]), 
        .A2(Red_SubCellInst_LFInst_13_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_13_LFInst_2_U2 ( .A(PermutationOutput[52]), 
        .ZN(Red_SubCellInst_LFInst_13_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_2_U1 ( .A1(PermutationOutput[53]), 
        .A2(PermutationOutput[52]), .ZN(Red_SubCellInst_LFInst_13_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U3 ( .A(PermutationOutput[57]), 
        .B(Red_SubCellInst_LFInst_14_LFInst_0_n2), .Z(Red_Feedback[42]) );
  OAI21_X1 Red_SubCellInst_LFInst_14_LFInst_0_U2 ( .B1(PermutationOutput[59]), 
        .B2(PermutationOutput[58]), .A(Red_SubCellInst_LFInst_14_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U1 ( .A1(PermutationOutput[59]), 
        .A2(PermutationOutput[56]), .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_14_LFInst_1_U5 ( .A1(PermutationOutput[56]), 
        .A2(Red_SubCellInst_LFInst_14_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_14_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_14_LFInst_1_n2), .ZN(Red_Feedback[43]) );
  OAI21_X1 Red_SubCellInst_LFInst_14_LFInst_1_U4 ( .B1(PermutationOutput[57]), 
        .B2(PermutationOutput[58]), .A(PermutationOutput[56]), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_14_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_14_LFInst_1_n2), .B(PermutationOutput[58]), .Z(
        Red_SubCellInst_LFInst_14_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_14_LFInst_1_U2 ( .A1(PermutationOutput[59]), 
        .A2(Red_SubCellInst_LFInst_14_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_14_LFInst_1_U1 ( .A(PermutationOutput[57]), 
        .ZN(Red_SubCellInst_LFInst_14_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_14_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_14_LFInst_2_n6), .B2(PermutationOutput[58]), 
        .C1(Red_SubCellInst_LFInst_14_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_14_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_14_LFInst_2_n3), .ZN(Red_Feedback[44]) );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_14_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U5 ( .A1(PermutationOutput[57]), 
        .A2(Red_SubCellInst_LFInst_14_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_14_LFInst_2_U4 ( .A(PermutationOutput[59]), 
        .ZN(Red_SubCellInst_LFInst_14_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U3 ( .A1(PermutationOutput[58]), 
        .A2(Red_SubCellInst_LFInst_14_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_14_LFInst_2_U2 ( .A(PermutationOutput[56]), 
        .ZN(Red_SubCellInst_LFInst_14_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_2_U1 ( .A1(PermutationOutput[57]), 
        .A2(PermutationOutput[56]), .ZN(Red_SubCellInst_LFInst_14_LFInst_2_n6)
         );
  XOR2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U3 ( .A(PermutationOutput[61]), 
        .B(Red_SubCellInst_LFInst_15_LFInst_0_n2), .Z(Red_Feedback[45]) );
  OAI21_X1 Red_SubCellInst_LFInst_15_LFInst_0_U2 ( .B1(PermutationOutput[63]), 
        .B2(PermutationOutput[62]), .A(Red_SubCellInst_LFInst_15_LFInst_0_n1), 
        .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U1 ( .A1(PermutationOutput[63]), 
        .A2(PermutationOutput[60]), .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n1)
         );
  OAI22_X1 Red_SubCellInst_LFInst_15_LFInst_1_U5 ( .A1(PermutationOutput[60]), 
        .A2(Red_SubCellInst_LFInst_15_LFInst_1_n4), .B1(
        Red_SubCellInst_LFInst_15_LFInst_1_n3), .B2(
        Red_SubCellInst_LFInst_15_LFInst_1_n2), .ZN(Red_Feedback[46]) );
  OAI21_X1 Red_SubCellInst_LFInst_15_LFInst_1_U4 ( .B1(PermutationOutput[61]), 
        .B2(PermutationOutput[62]), .A(PermutationOutput[60]), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_1_n3) );
  XOR2_X1 Red_SubCellInst_LFInst_15_LFInst_1_U3 ( .A(
        Red_SubCellInst_LFInst_15_LFInst_1_n2), .B(PermutationOutput[62]), .Z(
        Red_SubCellInst_LFInst_15_LFInst_1_n4) );
  NOR2_X1 Red_SubCellInst_LFInst_15_LFInst_1_U2 ( .A1(PermutationOutput[63]), 
        .A2(Red_SubCellInst_LFInst_15_LFInst_1_n1), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_1_n2) );
  INV_X1 Red_SubCellInst_LFInst_15_LFInst_1_U1 ( .A(PermutationOutput[61]), 
        .ZN(Red_SubCellInst_LFInst_15_LFInst_1_n1) );
  OAI221_X1 Red_SubCellInst_LFInst_15_LFInst_2_U7 ( .B1(
        Red_SubCellInst_LFInst_15_LFInst_2_n6), .B2(PermutationOutput[62]), 
        .C1(Red_SubCellInst_LFInst_15_LFInst_2_n5), .C2(
        Red_SubCellInst_LFInst_15_LFInst_2_n4), .A(
        Red_SubCellInst_LFInst_15_LFInst_2_n3), .ZN(Red_Feedback[47]) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U6 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_2_n5), .A2(
        Red_SubCellInst_LFInst_15_LFInst_2_n4), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_2_n3) );
  NOR2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U5 ( .A1(PermutationOutput[61]), 
        .A2(Red_SubCellInst_LFInst_15_LFInst_2_n2), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_2_n4) );
  INV_X1 Red_SubCellInst_LFInst_15_LFInst_2_U4 ( .A(PermutationOutput[63]), 
        .ZN(Red_SubCellInst_LFInst_15_LFInst_2_n2) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U3 ( .A1(PermutationOutput[62]), 
        .A2(Red_SubCellInst_LFInst_15_LFInst_2_n1), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_2_n5) );
  INV_X1 Red_SubCellInst_LFInst_15_LFInst_2_U2 ( .A(PermutationOutput[60]), 
        .ZN(Red_SubCellInst_LFInst_15_LFInst_2_n1) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_2_U1 ( .A1(PermutationOutput[61]), 
        .A2(PermutationOutput[60]), .ZN(Red_SubCellInst_LFInst_15_LFInst_2_n6)
         );
  BUF_X1 KeyMUX_U3 ( .A(selects[0]), .Z(KeyMUX_n2) );
  BUF_X1 KeyMUX_U2 ( .A(selects[0]), .Z(KeyMUX_n1) );
  BUF_X1 KeyMUX_U1 ( .A(selects[0]), .Z(KeyMUX_n3) );
  MUX2_X1 KeyMUX_MUXInst_0_U1 ( .A(Key[64]), .B(Key[0]), .S(KeyMUX_n1), .Z(
        SelectedKey[0]) );
  MUX2_X1 KeyMUX_MUXInst_1_U1 ( .A(Key[65]), .B(Key[1]), .S(KeyMUX_n2), .Z(
        SelectedKey[1]) );
  MUX2_X1 KeyMUX_MUXInst_2_U1 ( .A(Key[66]), .B(Key[2]), .S(KeyMUX_n2), .Z(
        SelectedKey[2]) );
  MUX2_X1 KeyMUX_MUXInst_3_U1 ( .A(Key[67]), .B(Key[3]), .S(KeyMUX_n2), .Z(
        SelectedKey[3]) );
  MUX2_X1 KeyMUX_MUXInst_4_U1 ( .A(Key[68]), .B(Key[4]), .S(KeyMUX_n2), .Z(
        SelectedKey[4]) );
  MUX2_X1 KeyMUX_MUXInst_5_U1 ( .A(Key[69]), .B(Key[5]), .S(selects[0]), .Z(
        SelectedKey[5]) );
  MUX2_X1 KeyMUX_MUXInst_6_U1 ( .A(Key[70]), .B(Key[6]), .S(KeyMUX_n2), .Z(
        SelectedKey[6]) );
  MUX2_X1 KeyMUX_MUXInst_7_U1 ( .A(Key[71]), .B(Key[7]), .S(selects[0]), .Z(
        SelectedKey[7]) );
  MUX2_X1 KeyMUX_MUXInst_8_U1 ( .A(Key[72]), .B(Key[8]), .S(KeyMUX_n2), .Z(
        SelectedKey[8]) );
  MUX2_X1 KeyMUX_MUXInst_9_U1 ( .A(Key[73]), .B(Key[9]), .S(selects[0]), .Z(
        SelectedKey[9]) );
  MUX2_X1 KeyMUX_MUXInst_10_U1 ( .A(Key[74]), .B(Key[10]), .S(selects[0]), .Z(
        SelectedKey[10]) );
  MUX2_X1 KeyMUX_MUXInst_11_U1 ( .A(Key[75]), .B(Key[11]), .S(KeyMUX_n1), .Z(
        SelectedKey[11]) );
  MUX2_X1 KeyMUX_MUXInst_12_U1 ( .A(Key[76]), .B(Key[12]), .S(selects[0]), .Z(
        SelectedKey[12]) );
  MUX2_X1 KeyMUX_MUXInst_13_U1 ( .A(Key[77]), .B(Key[13]), .S(selects[0]), .Z(
        SelectedKey[13]) );
  MUX2_X1 KeyMUX_MUXInst_14_U1 ( .A(Key[78]), .B(Key[14]), .S(selects[0]), .Z(
        SelectedKey[14]) );
  MUX2_X1 KeyMUX_MUXInst_15_U1 ( .A(Key[79]), .B(Key[15]), .S(selects[0]), .Z(
        SelectedKey[15]) );
  MUX2_X1 KeyMUX_MUXInst_16_U1 ( .A(Key[80]), .B(Key[16]), .S(selects[0]), .Z(
        SelectedKey[16]) );
  MUX2_X1 KeyMUX_MUXInst_17_U1 ( .A(Key[81]), .B(Key[17]), .S(KeyMUX_n2), .Z(
        SelectedKey[17]) );
  MUX2_X1 KeyMUX_MUXInst_18_U1 ( .A(Key[82]), .B(Key[18]), .S(KeyMUX_n3), .Z(
        SelectedKey[18]) );
  MUX2_X1 KeyMUX_MUXInst_19_U1 ( .A(Key[83]), .B(Key[19]), .S(KeyMUX_n3), .Z(
        SelectedKey[19]) );
  MUX2_X1 KeyMUX_MUXInst_20_U1 ( .A(Key[84]), .B(Key[20]), .S(KeyMUX_n1), .Z(
        SelectedKey[20]) );
  MUX2_X1 KeyMUX_MUXInst_21_U1 ( .A(Key[85]), .B(Key[21]), .S(KeyMUX_n3), .Z(
        SelectedKey[21]) );
  MUX2_X1 KeyMUX_MUXInst_22_U1 ( .A(Key[86]), .B(Key[22]), .S(KeyMUX_n3), .Z(
        SelectedKey[22]) );
  MUX2_X1 KeyMUX_MUXInst_23_U1 ( .A(Key[87]), .B(Key[23]), .S(KeyMUX_n2), .Z(
        SelectedKey[23]) );
  MUX2_X1 KeyMUX_MUXInst_24_U1 ( .A(Key[88]), .B(Key[24]), .S(KeyMUX_n3), .Z(
        SelectedKey[24]) );
  MUX2_X1 KeyMUX_MUXInst_25_U1 ( .A(Key[89]), .B(Key[25]), .S(KeyMUX_n3), .Z(
        SelectedKey[25]) );
  MUX2_X1 KeyMUX_MUXInst_26_U1 ( .A(Key[90]), .B(Key[26]), .S(KeyMUX_n3), .Z(
        SelectedKey[26]) );
  MUX2_X1 KeyMUX_MUXInst_27_U1 ( .A(Key[91]), .B(Key[27]), .S(KeyMUX_n3), .Z(
        SelectedKey[27]) );
  MUX2_X1 KeyMUX_MUXInst_28_U1 ( .A(Key[92]), .B(Key[28]), .S(KeyMUX_n3), .Z(
        SelectedKey[28]) );
  MUX2_X1 KeyMUX_MUXInst_29_U1 ( .A(Key[93]), .B(Key[29]), .S(KeyMUX_n3), .Z(
        SelectedKey[29]) );
  MUX2_X1 KeyMUX_MUXInst_30_U1 ( .A(Key[94]), .B(Key[30]), .S(KeyMUX_n3), .Z(
        SelectedKey[30]) );
  MUX2_X1 KeyMUX_MUXInst_31_U1 ( .A(Key[95]), .B(Key[31]), .S(KeyMUX_n3), .Z(
        SelectedKey[31]) );
  MUX2_X1 KeyMUX_MUXInst_32_U1 ( .A(Key[96]), .B(Key[32]), .S(KeyMUX_n3), .Z(
        SelectedKey[32]) );
  MUX2_X1 KeyMUX_MUXInst_33_U1 ( .A(Key[97]), .B(Key[33]), .S(KeyMUX_n3), .Z(
        SelectedKey[33]) );
  MUX2_X1 KeyMUX_MUXInst_34_U1 ( .A(Key[98]), .B(Key[34]), .S(KeyMUX_n3), .Z(
        SelectedKey[34]) );
  MUX2_X1 KeyMUX_MUXInst_35_U1 ( .A(Key[99]), .B(Key[35]), .S(KeyMUX_n3), .Z(
        SelectedKey[35]) );
  MUX2_X1 KeyMUX_MUXInst_36_U1 ( .A(Key[100]), .B(Key[36]), .S(KeyMUX_n1), .Z(
        SelectedKey[36]) );
  MUX2_X1 KeyMUX_MUXInst_37_U1 ( .A(Key[101]), .B(Key[37]), .S(KeyMUX_n1), .Z(
        SelectedKey[37]) );
  MUX2_X1 KeyMUX_MUXInst_38_U1 ( .A(Key[102]), .B(Key[38]), .S(KeyMUX_n1), .Z(
        SelectedKey[38]) );
  MUX2_X1 KeyMUX_MUXInst_39_U1 ( .A(Key[103]), .B(Key[39]), .S(KeyMUX_n1), .Z(
        SelectedKey[39]) );
  MUX2_X1 KeyMUX_MUXInst_40_U1 ( .A(Key[104]), .B(Key[40]), .S(KeyMUX_n1), .Z(
        SelectedKey[40]) );
  MUX2_X1 KeyMUX_MUXInst_41_U1 ( .A(Key[105]), .B(Key[41]), .S(KeyMUX_n1), .Z(
        SelectedKey[41]) );
  MUX2_X1 KeyMUX_MUXInst_42_U1 ( .A(Key[106]), .B(Key[42]), .S(KeyMUX_n1), .Z(
        SelectedKey[42]) );
  MUX2_X1 KeyMUX_MUXInst_43_U1 ( .A(Key[107]), .B(Key[43]), .S(KeyMUX_n1), .Z(
        SelectedKey[43]) );
  MUX2_X1 KeyMUX_MUXInst_44_U1 ( .A(Key[108]), .B(Key[44]), .S(KeyMUX_n1), .Z(
        SelectedKey[44]) );
  MUX2_X1 KeyMUX_MUXInst_45_U1 ( .A(Key[109]), .B(Key[45]), .S(KeyMUX_n1), .Z(
        SelectedKey[45]) );
  MUX2_X1 KeyMUX_MUXInst_46_U1 ( .A(Key[110]), .B(Key[46]), .S(KeyMUX_n1), .Z(
        SelectedKey[46]) );
  MUX2_X1 KeyMUX_MUXInst_47_U1 ( .A(Key[111]), .B(Key[47]), .S(KeyMUX_n1), .Z(
        SelectedKey[47]) );
  MUX2_X1 KeyMUX_MUXInst_48_U1 ( .A(Key[112]), .B(Key[48]), .S(KeyMUX_n2), .Z(
        SelectedKey[48]) );
  MUX2_X1 KeyMUX_MUXInst_49_U1 ( .A(Key[113]), .B(Key[49]), .S(KeyMUX_n2), .Z(
        SelectedKey[49]) );
  MUX2_X1 KeyMUX_MUXInst_50_U1 ( .A(Key[114]), .B(Key[50]), .S(KeyMUX_n2), .Z(
        SelectedKey[50]) );
  MUX2_X1 KeyMUX_MUXInst_51_U1 ( .A(Key[115]), .B(Key[51]), .S(KeyMUX_n2), .Z(
        SelectedKey[51]) );
  MUX2_X1 KeyMUX_MUXInst_52_U1 ( .A(Key[116]), .B(Key[52]), .S(KeyMUX_n2), .Z(
        SelectedKey[52]) );
  MUX2_X1 KeyMUX_MUXInst_53_U1 ( .A(Key[117]), .B(Key[53]), .S(KeyMUX_n2), .Z(
        SelectedKey[53]) );
  MUX2_X1 KeyMUX_MUXInst_54_U1 ( .A(Key[118]), .B(Key[54]), .S(KeyMUX_n2), .Z(
        SelectedKey[54]) );
  MUX2_X1 KeyMUX_MUXInst_55_U1 ( .A(Key[119]), .B(Key[55]), .S(KeyMUX_n2), .Z(
        SelectedKey[55]) );
  MUX2_X1 KeyMUX_MUXInst_56_U1 ( .A(Key[120]), .B(Key[56]), .S(KeyMUX_n2), .Z(
        SelectedKey[56]) );
  MUX2_X1 KeyMUX_MUXInst_57_U1 ( .A(Key[121]), .B(Key[57]), .S(KeyMUX_n2), .Z(
        SelectedKey[57]) );
  MUX2_X1 KeyMUX_MUXInst_58_U1 ( .A(Key[122]), .B(Key[58]), .S(KeyMUX_n2), .Z(
        SelectedKey[58]) );
  MUX2_X1 KeyMUX_MUXInst_59_U1 ( .A(Key[123]), .B(Key[59]), .S(KeyMUX_n2), .Z(
        SelectedKey[59]) );
  MUX2_X1 KeyMUX_MUXInst_60_U1 ( .A(Key[124]), .B(Key[60]), .S(KeyMUX_n3), .Z(
        SelectedKey[60]) );
  MUX2_X1 KeyMUX_MUXInst_61_U1 ( .A(Key[125]), .B(Key[61]), .S(KeyMUX_n3), .Z(
        SelectedKey[61]) );
  MUX2_X1 KeyMUX_MUXInst_62_U1 ( .A(Key[126]), .B(Key[62]), .S(KeyMUX_n3), .Z(
        SelectedKey[62]) );
  MUX2_X1 KeyMUX_MUXInst_63_U1 ( .A(Key[127]), .B(Key[63]), .S(KeyMUX_n3), .Z(
        SelectedKey[63]) );
  XNOR2_X1 Red_K0Inst_LFInst_0_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_0_LFInst_0_n1), .B(Key[66]), .ZN(Red_K0[0]) );
  XNOR2_X1 Red_K0Inst_LFInst_0_LFInst_0_U1 ( .A(Key[64]), .B(Key[65]), .ZN(
        Red_K0Inst_LFInst_0_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_0_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_0_LFInst_1_n1), .B(Key[67]), .ZN(Red_K0[1]) );
  XNOR2_X1 Red_K0Inst_LFInst_0_LFInst_1_U1 ( .A(Key[64]), .B(Key[65]), .ZN(
        Red_K0Inst_LFInst_0_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_0_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_0_LFInst_2_n1), .B(Key[67]), .ZN(Red_K0[2]) );
  XNOR2_X1 Red_K0Inst_LFInst_0_LFInst_2_U1 ( .A(Key[65]), .B(Key[66]), .ZN(
        Red_K0Inst_LFInst_0_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_1_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_1_LFInst_0_n1), .B(Key[70]), .ZN(Red_K0[3]) );
  XNOR2_X1 Red_K0Inst_LFInst_1_LFInst_0_U1 ( .A(Key[68]), .B(Key[69]), .ZN(
        Red_K0Inst_LFInst_1_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_1_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_1_LFInst_1_n1), .B(Key[71]), .ZN(Red_K0[4]) );
  XNOR2_X1 Red_K0Inst_LFInst_1_LFInst_1_U1 ( .A(Key[68]), .B(Key[69]), .ZN(
        Red_K0Inst_LFInst_1_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_1_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_1_LFInst_2_n1), .B(Key[71]), .ZN(Red_K0[5]) );
  XNOR2_X1 Red_K0Inst_LFInst_1_LFInst_2_U1 ( .A(Key[69]), .B(Key[70]), .ZN(
        Red_K0Inst_LFInst_1_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_2_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_2_LFInst_0_n1), .B(Key[74]), .ZN(Red_K0[6]) );
  XNOR2_X1 Red_K0Inst_LFInst_2_LFInst_0_U1 ( .A(Key[72]), .B(Key[73]), .ZN(
        Red_K0Inst_LFInst_2_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_2_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_2_LFInst_1_n1), .B(Key[75]), .ZN(Red_K0[7]) );
  XNOR2_X1 Red_K0Inst_LFInst_2_LFInst_1_U1 ( .A(Key[72]), .B(Key[73]), .ZN(
        Red_K0Inst_LFInst_2_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_2_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_2_LFInst_2_n1), .B(Key[75]), .ZN(Red_K0[8]) );
  XNOR2_X1 Red_K0Inst_LFInst_2_LFInst_2_U1 ( .A(Key[73]), .B(Key[74]), .ZN(
        Red_K0Inst_LFInst_2_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_3_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_3_LFInst_0_n1), .B(Key[78]), .ZN(Red_K0[9]) );
  XNOR2_X1 Red_K0Inst_LFInst_3_LFInst_0_U1 ( .A(Key[76]), .B(Key[77]), .ZN(
        Red_K0Inst_LFInst_3_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_3_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_3_LFInst_1_n1), .B(Key[79]), .ZN(Red_K0[10]) );
  XNOR2_X1 Red_K0Inst_LFInst_3_LFInst_1_U1 ( .A(Key[76]), .B(Key[77]), .ZN(
        Red_K0Inst_LFInst_3_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_3_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_3_LFInst_2_n1), .B(Key[79]), .ZN(Red_K0[11]) );
  XNOR2_X1 Red_K0Inst_LFInst_3_LFInst_2_U1 ( .A(Key[77]), .B(Key[78]), .ZN(
        Red_K0Inst_LFInst_3_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_4_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_4_LFInst_0_n1), .B(Key[82]), .ZN(Red_K0[12]) );
  XNOR2_X1 Red_K0Inst_LFInst_4_LFInst_0_U1 ( .A(Key[80]), .B(Key[81]), .ZN(
        Red_K0Inst_LFInst_4_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_4_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_4_LFInst_1_n1), .B(Key[83]), .ZN(Red_K0[13]) );
  XNOR2_X1 Red_K0Inst_LFInst_4_LFInst_1_U1 ( .A(Key[80]), .B(Key[81]), .ZN(
        Red_K0Inst_LFInst_4_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_4_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_4_LFInst_2_n1), .B(Key[83]), .ZN(Red_K0[14]) );
  XNOR2_X1 Red_K0Inst_LFInst_4_LFInst_2_U1 ( .A(Key[81]), .B(Key[82]), .ZN(
        Red_K0Inst_LFInst_4_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_5_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_5_LFInst_0_n1), .B(Key[86]), .ZN(Red_K0[15]) );
  XNOR2_X1 Red_K0Inst_LFInst_5_LFInst_0_U1 ( .A(Key[84]), .B(Key[85]), .ZN(
        Red_K0Inst_LFInst_5_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_5_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_5_LFInst_1_n1), .B(Key[87]), .ZN(Red_K0[16]) );
  XNOR2_X1 Red_K0Inst_LFInst_5_LFInst_1_U1 ( .A(Key[84]), .B(Key[85]), .ZN(
        Red_K0Inst_LFInst_5_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_5_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_5_LFInst_2_n1), .B(Key[87]), .ZN(Red_K0[17]) );
  XNOR2_X1 Red_K0Inst_LFInst_5_LFInst_2_U1 ( .A(Key[85]), .B(Key[86]), .ZN(
        Red_K0Inst_LFInst_5_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_6_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_6_LFInst_0_n1), .B(Key[90]), .ZN(Red_K0[18]) );
  XNOR2_X1 Red_K0Inst_LFInst_6_LFInst_0_U1 ( .A(Key[88]), .B(Key[89]), .ZN(
        Red_K0Inst_LFInst_6_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_6_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_6_LFInst_1_n1), .B(Key[91]), .ZN(Red_K0[19]) );
  XNOR2_X1 Red_K0Inst_LFInst_6_LFInst_1_U1 ( .A(Key[88]), .B(Key[89]), .ZN(
        Red_K0Inst_LFInst_6_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_6_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_6_LFInst_2_n1), .B(Key[91]), .ZN(Red_K0[20]) );
  XNOR2_X1 Red_K0Inst_LFInst_6_LFInst_2_U1 ( .A(Key[89]), .B(Key[90]), .ZN(
        Red_K0Inst_LFInst_6_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_7_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_7_LFInst_0_n1), .B(Key[94]), .ZN(Red_K0[21]) );
  XNOR2_X1 Red_K0Inst_LFInst_7_LFInst_0_U1 ( .A(Key[92]), .B(Key[93]), .ZN(
        Red_K0Inst_LFInst_7_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_7_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_7_LFInst_1_n1), .B(Key[95]), .ZN(Red_K0[22]) );
  XNOR2_X1 Red_K0Inst_LFInst_7_LFInst_1_U1 ( .A(Key[92]), .B(Key[93]), .ZN(
        Red_K0Inst_LFInst_7_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_7_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_7_LFInst_2_n1), .B(Key[95]), .ZN(Red_K0[23]) );
  XNOR2_X1 Red_K0Inst_LFInst_7_LFInst_2_U1 ( .A(Key[93]), .B(Key[94]), .ZN(
        Red_K0Inst_LFInst_7_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_8_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_8_LFInst_0_n1), .B(Key[98]), .ZN(Red_K0[24]) );
  XNOR2_X1 Red_K0Inst_LFInst_8_LFInst_0_U1 ( .A(Key[96]), .B(Key[97]), .ZN(
        Red_K0Inst_LFInst_8_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_8_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_8_LFInst_1_n1), .B(Key[99]), .ZN(Red_K0[25]) );
  XNOR2_X1 Red_K0Inst_LFInst_8_LFInst_1_U1 ( .A(Key[96]), .B(Key[97]), .ZN(
        Red_K0Inst_LFInst_8_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_8_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_8_LFInst_2_n1), .B(Key[99]), .ZN(Red_K0[26]) );
  XNOR2_X1 Red_K0Inst_LFInst_8_LFInst_2_U1 ( .A(Key[97]), .B(Key[98]), .ZN(
        Red_K0Inst_LFInst_8_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_9_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_9_LFInst_0_n1), .B(Key[102]), .ZN(Red_K0[27]) );
  XNOR2_X1 Red_K0Inst_LFInst_9_LFInst_0_U1 ( .A(Key[100]), .B(Key[101]), .ZN(
        Red_K0Inst_LFInst_9_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_9_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_9_LFInst_1_n1), .B(Key[103]), .ZN(Red_K0[28]) );
  XNOR2_X1 Red_K0Inst_LFInst_9_LFInst_1_U1 ( .A(Key[100]), .B(Key[101]), .ZN(
        Red_K0Inst_LFInst_9_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_9_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_9_LFInst_2_n1), .B(Key[103]), .ZN(Red_K0[29]) );
  XNOR2_X1 Red_K0Inst_LFInst_9_LFInst_2_U1 ( .A(Key[101]), .B(Key[102]), .ZN(
        Red_K0Inst_LFInst_9_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_10_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_10_LFInst_0_n1), .B(Key[106]), .ZN(Red_K0[30]) );
  XNOR2_X1 Red_K0Inst_LFInst_10_LFInst_0_U1 ( .A(Key[104]), .B(Key[105]), .ZN(
        Red_K0Inst_LFInst_10_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_10_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_10_LFInst_1_n1), .B(Key[107]), .ZN(Red_K0[31]) );
  XNOR2_X1 Red_K0Inst_LFInst_10_LFInst_1_U1 ( .A(Key[104]), .B(Key[105]), .ZN(
        Red_K0Inst_LFInst_10_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_10_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_10_LFInst_2_n1), .B(Key[107]), .ZN(Red_K0[32]) );
  XNOR2_X1 Red_K0Inst_LFInst_10_LFInst_2_U1 ( .A(Key[105]), .B(Key[106]), .ZN(
        Red_K0Inst_LFInst_10_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_11_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_11_LFInst_0_n1), .B(Key[110]), .ZN(Red_K0[33]) );
  XNOR2_X1 Red_K0Inst_LFInst_11_LFInst_0_U1 ( .A(Key[108]), .B(Key[109]), .ZN(
        Red_K0Inst_LFInst_11_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_11_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_11_LFInst_1_n1), .B(Key[111]), .ZN(Red_K0[34]) );
  XNOR2_X1 Red_K0Inst_LFInst_11_LFInst_1_U1 ( .A(Key[108]), .B(Key[109]), .ZN(
        Red_K0Inst_LFInst_11_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_11_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_11_LFInst_2_n1), .B(Key[111]), .ZN(Red_K0[35]) );
  XNOR2_X1 Red_K0Inst_LFInst_11_LFInst_2_U1 ( .A(Key[109]), .B(Key[110]), .ZN(
        Red_K0Inst_LFInst_11_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_12_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_12_LFInst_0_n1), .B(Key[114]), .ZN(Red_K0[36]) );
  XNOR2_X1 Red_K0Inst_LFInst_12_LFInst_0_U1 ( .A(Key[112]), .B(Key[113]), .ZN(
        Red_K0Inst_LFInst_12_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_12_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_12_LFInst_1_n1), .B(Key[115]), .ZN(Red_K0[37]) );
  XNOR2_X1 Red_K0Inst_LFInst_12_LFInst_1_U1 ( .A(Key[112]), .B(Key[113]), .ZN(
        Red_K0Inst_LFInst_12_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_12_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_12_LFInst_2_n1), .B(Key[115]), .ZN(Red_K0[38]) );
  XNOR2_X1 Red_K0Inst_LFInst_12_LFInst_2_U1 ( .A(Key[113]), .B(Key[114]), .ZN(
        Red_K0Inst_LFInst_12_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_13_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_13_LFInst_0_n1), .B(Key[118]), .ZN(Red_K0[39]) );
  XNOR2_X1 Red_K0Inst_LFInst_13_LFInst_0_U1 ( .A(Key[116]), .B(Key[117]), .ZN(
        Red_K0Inst_LFInst_13_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_13_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_13_LFInst_1_n1), .B(Key[119]), .ZN(Red_K0[40]) );
  XNOR2_X1 Red_K0Inst_LFInst_13_LFInst_1_U1 ( .A(Key[116]), .B(Key[117]), .ZN(
        Red_K0Inst_LFInst_13_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_13_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_13_LFInst_2_n1), .B(Key[119]), .ZN(Red_K0[41]) );
  XNOR2_X1 Red_K0Inst_LFInst_13_LFInst_2_U1 ( .A(Key[117]), .B(Key[118]), .ZN(
        Red_K0Inst_LFInst_13_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_14_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_14_LFInst_0_n1), .B(Key[122]), .ZN(Red_K0[42]) );
  XNOR2_X1 Red_K0Inst_LFInst_14_LFInst_0_U1 ( .A(Key[120]), .B(Key[121]), .ZN(
        Red_K0Inst_LFInst_14_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_14_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_14_LFInst_1_n1), .B(Key[123]), .ZN(Red_K0[43]) );
  XNOR2_X1 Red_K0Inst_LFInst_14_LFInst_1_U1 ( .A(Key[120]), .B(Key[121]), .ZN(
        Red_K0Inst_LFInst_14_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_14_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_14_LFInst_2_n1), .B(Key[123]), .ZN(Red_K0[44]) );
  XNOR2_X1 Red_K0Inst_LFInst_14_LFInst_2_U1 ( .A(Key[121]), .B(Key[122]), .ZN(
        Red_K0Inst_LFInst_14_LFInst_2_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_15_LFInst_0_U2 ( .A(
        Red_K0Inst_LFInst_15_LFInst_0_n1), .B(Key[126]), .ZN(Red_K0[45]) );
  XNOR2_X1 Red_K0Inst_LFInst_15_LFInst_0_U1 ( .A(Key[124]), .B(Key[125]), .ZN(
        Red_K0Inst_LFInst_15_LFInst_0_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_15_LFInst_1_U2 ( .A(
        Red_K0Inst_LFInst_15_LFInst_1_n1), .B(Key[127]), .ZN(Red_K0[46]) );
  XNOR2_X1 Red_K0Inst_LFInst_15_LFInst_1_U1 ( .A(Key[124]), .B(Key[125]), .ZN(
        Red_K0Inst_LFInst_15_LFInst_1_n1) );
  XNOR2_X1 Red_K0Inst_LFInst_15_LFInst_2_U2 ( .A(
        Red_K0Inst_LFInst_15_LFInst_2_n1), .B(Key[127]), .ZN(Red_K0[47]) );
  XNOR2_X1 Red_K0Inst_LFInst_15_LFInst_2_U1 ( .A(Key[125]), .B(Key[126]), .ZN(
        Red_K0Inst_LFInst_15_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_0_LFInst_0_n1), .B(Key[2]), .ZN(Red_K1[0]) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_0_U1 ( .A(Key[0]), .B(Key[1]), .ZN(
        Red_K1Inst_LFInst_0_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_0_LFInst_1_n1), .B(Key[3]), .ZN(Red_K1[1]) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_1_U1 ( .A(Key[0]), .B(Key[1]), .ZN(
        Red_K1Inst_LFInst_0_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_0_LFInst_2_n1), .B(Key[3]), .ZN(Red_K1[2]) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_2_U1 ( .A(Key[1]), .B(Key[2]), .ZN(
        Red_K1Inst_LFInst_0_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_1_LFInst_0_n1), .B(Key[6]), .ZN(Red_K1[3]) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_0_U1 ( .A(Key[4]), .B(Key[5]), .ZN(
        Red_K1Inst_LFInst_1_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_1_LFInst_1_n1), .B(Key[7]), .ZN(Red_K1[4]) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_1_U1 ( .A(Key[4]), .B(Key[5]), .ZN(
        Red_K1Inst_LFInst_1_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_1_LFInst_2_n1), .B(Key[7]), .ZN(Red_K1[5]) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_2_U1 ( .A(Key[5]), .B(Key[6]), .ZN(
        Red_K1Inst_LFInst_1_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_2_LFInst_0_n1), .B(Key[10]), .ZN(Red_K1[6]) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_0_U1 ( .A(Key[8]), .B(Key[9]), .ZN(
        Red_K1Inst_LFInst_2_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_2_LFInst_1_n1), .B(Key[11]), .ZN(Red_K1[7]) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_1_U1 ( .A(Key[8]), .B(Key[9]), .ZN(
        Red_K1Inst_LFInst_2_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_2_LFInst_2_n1), .B(Key[11]), .ZN(Red_K1[8]) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_2_U1 ( .A(Key[9]), .B(Key[10]), .ZN(
        Red_K1Inst_LFInst_2_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_3_LFInst_0_n1), .B(Key[14]), .ZN(Red_K1[9]) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_0_U1 ( .A(Key[12]), .B(Key[13]), .ZN(
        Red_K1Inst_LFInst_3_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_3_LFInst_1_n1), .B(Key[15]), .ZN(Red_K1[10]) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_1_U1 ( .A(Key[12]), .B(Key[13]), .ZN(
        Red_K1Inst_LFInst_3_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_3_LFInst_2_n1), .B(Key[15]), .ZN(Red_K1[11]) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_2_U1 ( .A(Key[13]), .B(Key[14]), .ZN(
        Red_K1Inst_LFInst_3_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_4_LFInst_0_n1), .B(Key[18]), .ZN(Red_K1[12]) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_0_U1 ( .A(Key[16]), .B(Key[17]), .ZN(
        Red_K1Inst_LFInst_4_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_4_LFInst_1_n1), .B(Key[19]), .ZN(Red_K1[13]) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_1_U1 ( .A(Key[16]), .B(Key[17]), .ZN(
        Red_K1Inst_LFInst_4_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_4_LFInst_2_n1), .B(Key[19]), .ZN(Red_K1[14]) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_2_U1 ( .A(Key[17]), .B(Key[18]), .ZN(
        Red_K1Inst_LFInst_4_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_5_LFInst_0_n1), .B(Key[22]), .ZN(Red_K1[15]) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_0_U1 ( .A(Key[20]), .B(Key[21]), .ZN(
        Red_K1Inst_LFInst_5_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_5_LFInst_1_n1), .B(Key[23]), .ZN(Red_K1[16]) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_1_U1 ( .A(Key[20]), .B(Key[21]), .ZN(
        Red_K1Inst_LFInst_5_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_5_LFInst_2_n1), .B(Key[23]), .ZN(Red_K1[17]) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_2_U1 ( .A(Key[21]), .B(Key[22]), .ZN(
        Red_K1Inst_LFInst_5_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_6_LFInst_0_n1), .B(Key[26]), .ZN(Red_K1[18]) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_0_U1 ( .A(Key[24]), .B(Key[25]), .ZN(
        Red_K1Inst_LFInst_6_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_6_LFInst_1_n1), .B(Key[27]), .ZN(Red_K1[19]) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_1_U1 ( .A(Key[24]), .B(Key[25]), .ZN(
        Red_K1Inst_LFInst_6_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_6_LFInst_2_n1), .B(Key[27]), .ZN(Red_K1[20]) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_2_U1 ( .A(Key[25]), .B(Key[26]), .ZN(
        Red_K1Inst_LFInst_6_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_7_LFInst_0_n1), .B(Key[30]), .ZN(Red_K1[21]) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_0_U1 ( .A(Key[28]), .B(Key[29]), .ZN(
        Red_K1Inst_LFInst_7_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_7_LFInst_1_n1), .B(Key[31]), .ZN(Red_K1[22]) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_1_U1 ( .A(Key[28]), .B(Key[29]), .ZN(
        Red_K1Inst_LFInst_7_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_7_LFInst_2_n1), .B(Key[31]), .ZN(Red_K1[23]) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_2_U1 ( .A(Key[29]), .B(Key[30]), .ZN(
        Red_K1Inst_LFInst_7_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_8_LFInst_0_n1), .B(Key[34]), .ZN(Red_K1[24]) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_0_U1 ( .A(Key[32]), .B(Key[33]), .ZN(
        Red_K1Inst_LFInst_8_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_8_LFInst_1_n1), .B(Key[35]), .ZN(Red_K1[25]) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_1_U1 ( .A(Key[32]), .B(Key[33]), .ZN(
        Red_K1Inst_LFInst_8_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_8_LFInst_2_n1), .B(Key[35]), .ZN(Red_K1[26]) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_2_U1 ( .A(Key[33]), .B(Key[34]), .ZN(
        Red_K1Inst_LFInst_8_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_9_LFInst_0_n1), .B(Key[38]), .ZN(Red_K1[27]) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_0_U1 ( .A(Key[36]), .B(Key[37]), .ZN(
        Red_K1Inst_LFInst_9_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_9_LFInst_1_n1), .B(Key[39]), .ZN(Red_K1[28]) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_1_U1 ( .A(Key[36]), .B(Key[37]), .ZN(
        Red_K1Inst_LFInst_9_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_9_LFInst_2_n1), .B(Key[39]), .ZN(Red_K1[29]) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_2_U1 ( .A(Key[37]), .B(Key[38]), .ZN(
        Red_K1Inst_LFInst_9_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_10_LFInst_0_n1), .B(Key[42]), .ZN(Red_K1[30]) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_0_U1 ( .A(Key[40]), .B(Key[41]), .ZN(
        Red_K1Inst_LFInst_10_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_10_LFInst_1_n1), .B(Key[43]), .ZN(Red_K1[31]) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_1_U1 ( .A(Key[40]), .B(Key[41]), .ZN(
        Red_K1Inst_LFInst_10_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_10_LFInst_2_n1), .B(Key[43]), .ZN(Red_K1[32]) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_2_U1 ( .A(Key[41]), .B(Key[42]), .ZN(
        Red_K1Inst_LFInst_10_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_11_LFInst_0_n1), .B(Key[46]), .ZN(Red_K1[33]) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_0_U1 ( .A(Key[44]), .B(Key[45]), .ZN(
        Red_K1Inst_LFInst_11_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_11_LFInst_1_n1), .B(Key[47]), .ZN(Red_K1[34]) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_1_U1 ( .A(Key[44]), .B(Key[45]), .ZN(
        Red_K1Inst_LFInst_11_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_11_LFInst_2_n1), .B(Key[47]), .ZN(Red_K1[35]) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_2_U1 ( .A(Key[45]), .B(Key[46]), .ZN(
        Red_K1Inst_LFInst_11_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_12_LFInst_0_n1), .B(Key[50]), .ZN(Red_K1[36]) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_0_U1 ( .A(Key[48]), .B(Key[49]), .ZN(
        Red_K1Inst_LFInst_12_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_12_LFInst_1_n1), .B(Key[51]), .ZN(Red_K1[37]) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_1_U1 ( .A(Key[48]), .B(Key[49]), .ZN(
        Red_K1Inst_LFInst_12_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_12_LFInst_2_n1), .B(Key[51]), .ZN(Red_K1[38]) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_2_U1 ( .A(Key[49]), .B(Key[50]), .ZN(
        Red_K1Inst_LFInst_12_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_13_LFInst_0_n1), .B(Key[54]), .ZN(Red_K1[39]) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_0_U1 ( .A(Key[52]), .B(Key[53]), .ZN(
        Red_K1Inst_LFInst_13_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_13_LFInst_1_n1), .B(Key[55]), .ZN(Red_K1[40]) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_1_U1 ( .A(Key[52]), .B(Key[53]), .ZN(
        Red_K1Inst_LFInst_13_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_13_LFInst_2_n1), .B(Key[55]), .ZN(Red_K1[41]) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_2_U1 ( .A(Key[53]), .B(Key[54]), .ZN(
        Red_K1Inst_LFInst_13_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_14_LFInst_0_n1), .B(Key[58]), .ZN(Red_K1[42]) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_0_U1 ( .A(Key[56]), .B(Key[57]), .ZN(
        Red_K1Inst_LFInst_14_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_14_LFInst_1_n1), .B(Key[59]), .ZN(Red_K1[43]) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_1_U1 ( .A(Key[56]), .B(Key[57]), .ZN(
        Red_K1Inst_LFInst_14_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_14_LFInst_2_n1), .B(Key[59]), .ZN(Red_K1[44]) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_2_U1 ( .A(Key[57]), .B(Key[58]), .ZN(
        Red_K1Inst_LFInst_14_LFInst_2_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_0_U2 ( .A(
        Red_K1Inst_LFInst_15_LFInst_0_n1), .B(Key[62]), .ZN(Red_K1[45]) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_0_U1 ( .A(Key[60]), .B(Key[61]), .ZN(
        Red_K1Inst_LFInst_15_LFInst_0_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_1_U2 ( .A(
        Red_K1Inst_LFInst_15_LFInst_1_n1), .B(Key[63]), .ZN(Red_K1[46]) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_1_U1 ( .A(Key[60]), .B(Key[61]), .ZN(
        Red_K1Inst_LFInst_15_LFInst_1_n1) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_2_U2 ( .A(
        Red_K1Inst_LFInst_15_LFInst_2_n1), .B(Key[63]), .ZN(Red_K1[47]) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_2_U1 ( .A(Key[61]), .B(Key[62]), .ZN(
        Red_K1Inst_LFInst_15_LFInst_2_n1) );
  BUF_X2 Red_KeyMUX_U6 ( .A(Red_sel_Key[0]), .Z(Red_KeyMUX_n1) );
  BUF_X1 Red_KeyMUX_U5 ( .A(Red_sel_Key[1]), .Z(Red_KeyMUX_n4) );
  BUF_X1 Red_KeyMUX_U4 ( .A(Red_sel_Key[2]), .Z(Red_KeyMUX_n6) );
  BUF_X1 Red_KeyMUX_U3 ( .A(Red_sel_Key[1]), .Z(Red_KeyMUX_n3) );
  BUF_X1 Red_KeyMUX_U2 ( .A(Red_sel_Key[2]), .Z(Red_KeyMUX_n5) );
  CLKBUF_X3 Red_KeyMUX_U1 ( .A(Red_sel_Key[0]), .Z(Red_KeyMUX_n2) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_0_MUXInst_0_0_U1 ( .A(Red_K0[0]), .B(1'b0), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_0_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_0_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[0]), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_0_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_0_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_0_S_1__0_), .B(Red_KeyMUX_MUX2to1Inst_0_S_1__1_), .S(Red_KeyMUX_n4), .Z(Red_KeyMUX_MUX2to1Inst_0_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_0_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_0_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[0]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_1_MUXInst_0_0_U1 ( .A(Red_K0[1]), .B(1'b0), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_1_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_1_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[1]), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_1_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_1_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_1_S_1__0_), .B(Red_KeyMUX_MUX2to1Inst_1_S_1__1_), .S(Red_KeyMUX_n4), .Z(Red_KeyMUX_MUX2to1Inst_1_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_1_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_1_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[1]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_2_MUXInst_0_0_U1 ( .A(Red_K0[2]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_2_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_2_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[2]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_2_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_2_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_2_S_1__0_), .B(Red_KeyMUX_MUX2to1Inst_2_S_1__1_), .S(Red_sel_Key[1]), .Z(Red_KeyMUX_MUX2to1Inst_2_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_2_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_2_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[2]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_3_MUXInst_0_0_U1 ( .A(Red_K0[3]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_3_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_3_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[3]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_3_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_3_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_3_S_1__0_), .B(Red_KeyMUX_MUX2to1Inst_3_S_1__1_), .S(Red_sel_Key[1]), .Z(Red_KeyMUX_MUX2to1Inst_3_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_3_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_3_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[3]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_4_MUXInst_0_0_U1 ( .A(Red_K0[4]), .B(1'b0), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_4_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_4_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[4]), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_4_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_4_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_4_S_1__0_), .B(Red_KeyMUX_MUX2to1Inst_4_S_1__1_), .S(Red_KeyMUX_n4), .Z(Red_KeyMUX_MUX2to1Inst_4_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_4_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_4_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[4]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_5_MUXInst_0_0_U1 ( .A(Red_K0[5]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_5_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_5_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[5]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_5_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_5_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_5_S_1__0_), .B(Red_KeyMUX_MUX2to1Inst_5_S_1__1_), .S(Red_KeyMUX_n4), .Z(Red_KeyMUX_MUX2to1Inst_5_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_5_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_5_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[5]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_6_MUXInst_0_0_U1 ( .A(Red_K0[6]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_6_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_6_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[6]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_6_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_6_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_6_S_1__0_), .B(Red_KeyMUX_MUX2to1Inst_6_S_1__1_), .S(Red_KeyMUX_n4), .Z(Red_KeyMUX_MUX2to1Inst_6_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_6_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_6_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[6]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_7_MUXInst_0_0_U1 ( .A(Red_K0[7]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_7_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_7_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[7]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_7_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_7_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_7_S_1__0_), .B(Red_KeyMUX_MUX2to1Inst_7_S_1__1_), .S(Red_KeyMUX_n4), .Z(Red_KeyMUX_MUX2to1Inst_7_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_7_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_7_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[7]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_8_MUXInst_0_0_U1 ( .A(Red_K0[8]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_8_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_8_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[8]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_8_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_8_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_8_S_1__0_), .B(Red_KeyMUX_MUX2to1Inst_8_S_1__1_), .S(Red_sel_Key[1]), .Z(Red_KeyMUX_MUX2to1Inst_8_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_8_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_8_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[8]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_9_MUXInst_0_0_U1 ( .A(Red_K0[9]), .B(1'b0), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_9_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_9_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[9]), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_9_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_9_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_9_S_1__0_), .B(Red_KeyMUX_MUX2to1Inst_9_S_1__1_), .S(Red_sel_Key[1]), .Z(Red_KeyMUX_MUX2to1Inst_9_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_9_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_9_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[9]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_10_MUXInst_0_0_U1 ( .A(Red_K0[10]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_10_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_10_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[10]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_10_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_10_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_10_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_10_S_1__1_), .S(Red_KeyMUX_n4), .Z(
        Red_KeyMUX_MUX2to1Inst_10_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_10_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_10_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[10]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_11_MUXInst_0_0_U1 ( .A(Red_K0[11]), .B(1'b0), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_11_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_11_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[11]), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_11_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_11_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_11_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_11_S_1__1_), .S(Red_KeyMUX_n4), .Z(
        Red_KeyMUX_MUX2to1Inst_11_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_11_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_11_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[11]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_12_MUXInst_0_0_U1 ( .A(Red_K0[12]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_12_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_12_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[12]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_12_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_12_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_12_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_12_S_1__1_), .S(Red_sel_Key[1]), .Z(
        Red_KeyMUX_MUX2to1Inst_12_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_12_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_12_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[12]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_13_MUXInst_0_0_U1 ( .A(Red_K0[13]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_13_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_13_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[13]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_13_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_13_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_13_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_13_S_1__1_), .S(Red_sel_Key[1]), .Z(
        Red_KeyMUX_MUX2to1Inst_13_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_13_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_13_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[13]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_14_MUXInst_0_0_U1 ( .A(Red_K0[14]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_14_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_14_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[14]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_14_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_14_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_14_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_14_S_1__1_), .S(Red_sel_Key[1]), .Z(
        Red_KeyMUX_MUX2to1Inst_14_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_14_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_14_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[14]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_15_MUXInst_0_0_U1 ( .A(Red_K0[15]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_15_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_15_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[15]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_15_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_15_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_15_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_15_S_1__1_), .S(Red_sel_Key[1]), .Z(
        Red_KeyMUX_MUX2to1Inst_15_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_15_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_15_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[15]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_16_MUXInst_0_0_U1 ( .A(Red_K0[16]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_16_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_16_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[16]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_16_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_16_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_16_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_16_S_1__1_), .S(Red_sel_Key[1]), .Z(
        Red_KeyMUX_MUX2to1Inst_16_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_16_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_16_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[16]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_17_MUXInst_0_0_U1 ( .A(Red_K0[17]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_17_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_17_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[17]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_17_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_17_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_17_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_17_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_17_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_17_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_17_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[17]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_18_MUXInst_0_0_U1 ( .A(Red_K0[18]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_18_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_18_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[18]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_18_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_18_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_18_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_18_S_1__1_), .S(Red_sel_Key[1]), .Z(
        Red_KeyMUX_MUX2to1Inst_18_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_18_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_18_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[18]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_19_MUXInst_0_0_U1 ( .A(Red_K0[19]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_19_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_19_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[19]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_19_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_19_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_19_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_19_S_1__1_), .S(Red_sel_Key[1]), .Z(
        Red_KeyMUX_MUX2to1Inst_19_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_19_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_19_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[19]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_20_MUXInst_0_0_U1 ( .A(Red_K0[20]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_20_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_20_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[20]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_20_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_20_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_20_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_20_S_1__1_), .S(Red_sel_Key[1]), .Z(
        Red_KeyMUX_MUX2to1Inst_20_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_20_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_20_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[20]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_21_MUXInst_0_0_U1 ( .A(Red_K0[21]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_21_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_21_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[21]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_21_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_21_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_21_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_21_S_1__1_), .S(Red_sel_Key[1]), .Z(
        Red_KeyMUX_MUX2to1Inst_21_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_21_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_21_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[21]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_22_MUXInst_0_0_U1 ( .A(Red_K0[22]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_22_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_22_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[22]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_22_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_22_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_22_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_22_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_22_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_22_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_22_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[22]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_23_MUXInst_0_0_U1 ( .A(Red_K0[23]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_23_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_23_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[23]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_23_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_23_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_23_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_23_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_23_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_23_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_23_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[23]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_24_MUXInst_0_0_U1 ( .A(Red_K0[24]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_24_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_24_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[24]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_24_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_24_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_24_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_24_S_1__1_), .S(Red_sel_Key[1]), .Z(
        Red_KeyMUX_MUX2to1Inst_24_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_24_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_24_S_2__0_), .B(1'b0), .S(Red_sel_Key[2]), .Z(
        Red_SelectedKey[24]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_25_MUXInst_0_0_U1 ( .A(Red_K0[25]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_25_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_25_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[25]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_25_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_25_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_25_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_25_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_25_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_25_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_25_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[25]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_26_MUXInst_0_0_U1 ( .A(Red_K0[26]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_26_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_26_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[26]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_26_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_26_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_26_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_26_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_26_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_26_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_26_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[26]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_27_MUXInst_0_0_U1 ( .A(Red_K0[27]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_27_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_27_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[27]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_27_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_27_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_27_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_27_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_27_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_27_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_27_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[27]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_28_MUXInst_0_0_U1 ( .A(Red_K0[28]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_28_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_28_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[28]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_28_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_28_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_28_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_28_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_28_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_28_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_28_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[28]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_29_MUXInst_0_0_U1 ( .A(Red_K0[29]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_29_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_29_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[29]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_29_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_29_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_29_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_29_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_29_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_29_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_29_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[29]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_30_MUXInst_0_0_U1 ( .A(Red_K0[30]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_30_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_30_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[30]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_30_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_30_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_30_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_30_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_30_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_30_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_30_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[30]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_31_MUXInst_0_0_U1 ( .A(Red_K0[31]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_31_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_31_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[31]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_31_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_31_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_31_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_31_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_31_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_31_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_31_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[31]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_32_MUXInst_0_0_U1 ( .A(Red_K0[32]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_32_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_32_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[32]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_32_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_32_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_32_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_32_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_32_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_32_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_32_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[32]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_33_MUXInst_0_0_U1 ( .A(Red_K0[33]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_33_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_33_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[33]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_33_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_33_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_33_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_33_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_33_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_33_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_33_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[33]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_34_MUXInst_0_0_U1 ( .A(Red_K0[34]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_34_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_34_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[34]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_34_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_34_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_34_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_34_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_34_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_34_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_34_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[34]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_35_MUXInst_0_0_U1 ( .A(Red_K0[35]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_35_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_35_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[35]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_35_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_35_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_35_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_35_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_35_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_35_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_35_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[35]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_36_MUXInst_0_0_U1 ( .A(Red_K0[36]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_36_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_36_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[36]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_36_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_36_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_36_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_36_S_1__1_), .S(Red_KeyMUX_n3), .Z(
        Red_KeyMUX_MUX2to1Inst_36_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_36_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_36_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n5), .Z(
        Red_SelectedKey[36]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_37_MUXInst_0_0_U1 ( .A(Red_K0[37]), .B(1'b0), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_37_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_37_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[37]), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_37_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_37_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_37_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_37_S_1__1_), .S(Red_KeyMUX_n4), .Z(
        Red_KeyMUX_MUX2to1Inst_37_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_37_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_37_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[37]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_38_MUXInst_0_0_U1 ( .A(Red_K0[38]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_38_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_38_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[38]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_38_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_38_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_38_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_38_S_1__1_), .S(Red_KeyMUX_n4), .Z(
        Red_KeyMUX_MUX2to1Inst_38_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_38_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_38_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[38]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_39_MUXInst_0_0_U1 ( .A(Red_K0[39]), .B(1'b0), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_39_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_39_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[39]), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_39_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_39_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_39_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_39_S_1__1_), .S(Red_KeyMUX_n4), .Z(
        Red_KeyMUX_MUX2to1Inst_39_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_39_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_39_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[39]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_40_MUXInst_0_0_U1 ( .A(Red_K0[40]), .B(1'b0), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_40_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_40_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[40]), 
        .S(Red_sel_Key[0]), .Z(Red_KeyMUX_MUX2to1Inst_40_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_40_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_40_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_40_S_1__1_), .S(Red_KeyMUX_n4), .Z(
        Red_KeyMUX_MUX2to1Inst_40_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_40_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_40_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[40]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_41_MUXInst_0_0_U1 ( .A(Red_K0[41]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_41_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_41_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[41]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_41_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_41_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_41_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_41_S_1__1_), .S(Red_KeyMUX_n4), .Z(
        Red_KeyMUX_MUX2to1Inst_41_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_41_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_41_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[41]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_42_MUXInst_0_0_U1 ( .A(Red_K0[42]), .B(1'b0), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_42_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_42_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[42]), 
        .S(Red_KeyMUX_n1), .Z(Red_KeyMUX_MUX2to1Inst_42_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_42_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_42_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_42_S_1__1_), .S(Red_KeyMUX_n4), .Z(
        Red_KeyMUX_MUX2to1Inst_42_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_42_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_42_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[42]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_43_MUXInst_0_0_U1 ( .A(Red_K0[43]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_43_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_43_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[43]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_43_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_43_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_43_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_43_S_1__1_), .S(Red_KeyMUX_n4), .Z(
        Red_KeyMUX_MUX2to1Inst_43_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_43_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_43_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[43]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_44_MUXInst_0_0_U1 ( .A(Red_K0[44]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_44_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_44_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[44]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_44_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_44_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_44_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_44_S_1__1_), .S(Red_KeyMUX_n4), .Z(
        Red_KeyMUX_MUX2to1Inst_44_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_44_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_44_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[44]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_45_MUXInst_0_0_U1 ( .A(Red_K0[45]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_45_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_45_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[45]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_45_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_45_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_45_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_45_S_1__1_), .S(Red_KeyMUX_n4), .Z(
        Red_KeyMUX_MUX2to1Inst_45_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_45_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_45_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[45]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_46_MUXInst_0_0_U1 ( .A(Red_K0[46]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_46_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_46_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[46]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_46_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_46_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_46_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_46_S_1__1_), .S(Red_KeyMUX_n4), .Z(
        Red_KeyMUX_MUX2to1Inst_46_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_46_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_46_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[46]) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_47_MUXInst_0_0_U1 ( .A(Red_K0[47]), .B(1'b0), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_47_S_1__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_47_MUXInst_0_1_U1 ( .A(1'b0), .B(Red_K1[47]), 
        .S(Red_KeyMUX_n2), .Z(Red_KeyMUX_MUX2to1Inst_47_S_1__1_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_47_MUXInst_1_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_47_S_1__0_), .B(
        Red_KeyMUX_MUX2to1Inst_47_S_1__1_), .S(Red_KeyMUX_n4), .Z(
        Red_KeyMUX_MUX2to1Inst_47_S_2__0_) );
  MUX2_X1 Red_KeyMUX_MUX2to1Inst_47_MUXInst_2_0_U1 ( .A(
        Red_KeyMUX_MUX2to1Inst_47_S_2__0_), .B(1'b0), .S(Red_KeyMUX_n6), .Z(
        Red_SelectedKey[47]) );
  MUX2_X1 FSMMUX_MUXInst_0_U1 ( .A(FSMReg[0]), .B(1'b1), .S(rst), .Z(
        RoundConstant_0) );
  MUX2_X1 FSMMUX_MUXInst_1_U1 ( .A(FSMReg[1]), .B(1'b0), .S(rst), .Z(
        FSMUpdate[0]) );
  MUX2_X1 FSMMUX_MUXInst_2_U1 ( .A(FSMReg[2]), .B(1'b0), .S(rst), .Z(
        FSMUpdate[1]) );
  MUX2_X1 FSMMUX_MUXInst_3_U1 ( .A(FSMReg[3]), .B(1'b1), .S(rst), .Z(
        RoundConstant_4_) );
  MUX2_X1 FSMMUX_MUXInst_4_U1 ( .A(FSMReg[4]), .B(1'b0), .S(rst), .Z(
        FSMUpdate[3]) );
  MUX2_X1 FSMMUX_MUXInst_5_U1 ( .A(FSMReg[5]), .B(1'b0), .S(rst), .Z(
        FSMUpdate[4]) );
  MUX2_X1 FSMMUX_MUXInst_6_U1 ( .A(FSMReg[6]), .B(1'b0), .S(rst), .Z(
        FSMUpdate[5]) );
  XOR2_X1 FSMUpdateInst_StateUpdateBitInst_2_U1 ( .A(RoundConstant_0), .B(
        FSMUpdate[0]), .Z(FSMUpdate[2]) );
  XOR2_X1 FSMUpdateInst_StateUpdateBitInst_6_U1 ( .A(RoundConstant_4_), .B(
        FSMUpdate[3]), .Z(FSMUpdate[6]) );
  DFF_X1 FSMRegInst_s_current_state_reg_0_ ( .D(FSMUpdate[0]), .CK(clk), .Q(
        FSMReg[0]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_1_ ( .D(FSMUpdate[1]), .CK(clk), .Q(
        FSMReg[1]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_2_ ( .D(FSMUpdate[2]), .CK(clk), .Q(
        FSMReg[2]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_3_ ( .D(FSMUpdate[3]), .CK(clk), .Q(
        FSMReg[3]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_4_ ( .D(FSMUpdate[4]), .CK(clk), .Q(
        FSMReg[4]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_5_ ( .D(FSMUpdate[5]), .CK(clk), .Q(
        FSMReg[5]), .QN() );
  DFF_X1 FSMRegInst_s_current_state_reg_6_ ( .D(FSMUpdate[6]), .CK(clk), .Q(
        FSMReg[6]), .QN() );
  NOR4_X1 FSMSignals_doneInst_U2 ( .A1(RoundConstant_0), .A2(RoundConstant_4_), 
        .A3(FSMUpdate[3]), .A4(FSMUpdate[5]), .ZN(FSMSignals_doneInst_n1) );
  AND4_X1 FSMSignals_doneInst_U1 ( .A1(FSMUpdate[0]), .A2(FSMUpdate[1]), .A3(
        FSMUpdate[4]), .A4(FSMSignals_doneInst_n1), .ZN(done) );
  MUX2_X1 selectsMUX_MUXInst_0_U1 ( .A(selectsReg[0]), .B(1'b0), .S(rst), .Z(
        selects[0]) );
  MUX2_X1 selectsMUX_MUXInst_1_U1 ( .A(selectsReg[1]), .B(1'b0), .S(rst), .Z(
        selects[1]) );
  INV_X1 selectsUpdateInst_selectsUpdateBitInst_0_U1 ( .A(selects[0]), .ZN(
        selectsNext[0]) );
  XOR2_X1 selectsUpdateInst_selectsUpdateBitInst_1_U1 ( .A(selects[0]), .B(
        selects[1]), .Z(selectsNext[1]) );
  DFF_X1 selectsRegInst_s_current_state_reg_0_ ( .D(selectsNext[0]), .CK(clk), 
        .Q(selectsReg[0]), .QN() );
  DFF_X1 selectsRegInst_s_current_state_reg_1_ ( .D(selectsNext[1]), .CK(clk), 
        .Q(selectsReg[1]), .QN() );
  MUX2_X1 Red_FSMMUX_MUXInst_0_U1 ( .A(Red_FSMReg[0]), .B(1'b1), .S(rst), .Z(
        Red_RoundConstant[0]) );
  MUX2_X1 Red_FSMMUX_MUXInst_1_U1 ( .A(Red_FSMReg[1]), .B(1'b1), .S(rst), .Z(
        Red_RoundConstant[1]) );
  MUX2_X1 Red_FSMMUX_MUXInst_2_U1 ( .A(Red_FSMReg[2]), .B(1'b0), .S(rst), .Z(
        Red_RoundConstant[2]) );
  MUX2_X1 Red_FSMMUX_MUXInst_3_U1 ( .A(Red_FSMReg[3]), .B(1'b1), .S(rst), .Z(
        Red_RoundConstant[3]) );
  MUX2_X1 Red_FSMMUX_MUXInst_4_U1 ( .A(Red_FSMReg[4]), .B(1'b1), .S(rst), .Z(
        Red_RoundConstant[4]) );
  MUX2_X1 Red_FSMMUX_MUXInst_5_U1 ( .A(Red_FSMReg[5]), .B(1'b0), .S(rst), .Z(
        Red_RoundConstant[5]) );
  XOR2_X1 Red_FSMUpdateInst_Red_StateUpdateBitInst_0_U2 ( .A(RoundConstant_0), 
        .B(FSMUpdate[1]), .Z(Red_FSMUpdate[0]) );
  XOR2_X1 Red_FSMUpdateInst_Red_StateUpdateBitInst_1_U2 ( .A(FSMUpdate[0]), 
        .B(FSMUpdate[1]), .Z(Red_FSMUpdate[1]) );
  XNOR2_X1 Red_FSMUpdateInst_Red_StateUpdateBitInst_2_U3 ( .A(
        Red_FSMUpdateInst_Red_StateUpdateBitInst_2_n1), .B(FSMUpdate[1]), .ZN(
        Red_FSMUpdate[2]) );
  XNOR2_X1 Red_FSMUpdateInst_Red_StateUpdateBitInst_2_U2 ( .A(RoundConstant_0), 
        .B(FSMUpdate[0]), .ZN(Red_FSMUpdateInst_Red_StateUpdateBitInst_2_n1)
         );
  XNOR2_X1 Red_FSMUpdateInst_Red_StateUpdateBitInst_3_U2 ( .A(
        Red_FSMUpdateInst_Red_StateUpdateBitInst_3_n1), .B(FSMUpdate[5]), .ZN(
        Red_FSMUpdate[3]) );
  XNOR2_X1 Red_FSMUpdateInst_Red_StateUpdateBitInst_3_U1 ( .A(FSMUpdate[3]), 
        .B(FSMUpdate[4]), .ZN(Red_FSMUpdateInst_Red_StateUpdateBitInst_3_n1)
         );
  XOR2_X1 Red_FSMUpdateInst_Red_StateUpdateBitInst_4_U1 ( .A(RoundConstant_4_), 
        .B(FSMUpdate[4]), .Z(Red_FSMUpdate[4]) );
  XNOR2_X1 Red_FSMUpdateInst_Red_StateUpdateBitInst_5_U3 ( .A(
        Red_FSMUpdateInst_Red_StateUpdateBitInst_5_n2), .B(
        Red_FSMUpdateInst_Red_StateUpdateBitInst_5_n1), .ZN(Red_FSMUpdate[5])
         );
  XNOR2_X1 Red_FSMUpdateInst_Red_StateUpdateBitInst_5_U2 ( .A(FSMUpdate[4]), 
        .B(FSMUpdate[5]), .ZN(Red_FSMUpdateInst_Red_StateUpdateBitInst_5_n1)
         );
  XOR2_X1 Red_FSMUpdateInst_Red_StateUpdateBitInst_5_U1 ( .A(RoundConstant_4_), 
        .B(FSMUpdate[3]), .Z(Red_FSMUpdateInst_Red_StateUpdateBitInst_5_n2) );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_0_ ( .D(Red_FSMUpdate[0]), .CK(clk), .Q(Red_FSMReg[0]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_1_ ( .D(Red_FSMUpdate[1]), .CK(clk), .Q(Red_FSMReg[1]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_2_ ( .D(Red_FSMUpdate[2]), .CK(clk), .Q(Red_FSMReg[2]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_3_ ( .D(Red_FSMUpdate[3]), .CK(clk), .Q(Red_FSMReg[3]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_4_ ( .D(Red_FSMUpdate[4]), .CK(clk), .Q(Red_FSMReg[4]), .QN() );
  DFF_X1 Red_FSMRegInst_s_current_state_reg_5_ ( .D(Red_FSMUpdate[5]), .CK(clk), .Q(Red_FSMReg[5]), .QN() );
  AND4_X1 Red_FSMSignals_doneInst_Red_FSMSignals_doneBitInst_0_U3 ( .A1(
        FSMUpdate[0]), .A2(FSMUpdate[1]), .A3(FSMUpdate[4]), .A4(
        Red_FSMSignals_doneInst_Red_FSMSignals_doneBitInst_0_n1), .ZN(
        Red_done[0]) );
  NOR4_X1 Red_FSMSignals_doneInst_Red_FSMSignals_doneBitInst_0_U2 ( .A1(
        RoundConstant_0), .A2(RoundConstant_4_), .A3(FSMUpdate[3]), .A4(
        FSMUpdate[5]), .ZN(
        Red_FSMSignals_doneInst_Red_FSMSignals_doneBitInst_0_n1) );
  AND4_X1 Red_FSMSignals_doneInst_Red_FSMSignals_doneBitInst_1_U3 ( .A1(
        FSMUpdate[0]), .A2(FSMUpdate[1]), .A3(FSMUpdate[4]), .A4(
        Red_FSMSignals_doneInst_Red_FSMSignals_doneBitInst_1_n1), .ZN(
        Red_done[1]) );
  NOR4_X1 Red_FSMSignals_doneInst_Red_FSMSignals_doneBitInst_1_U2 ( .A1(
        RoundConstant_0), .A2(RoundConstant_4_), .A3(FSMUpdate[3]), .A4(
        FSMUpdate[5]), .ZN(
        Red_FSMSignals_doneInst_Red_FSMSignals_doneBitInst_1_n1) );
  MUX2_X1 Red_selectsMUX_MUXInst_0_U1 ( .A(Red_selectsReg[0]), .B(1'b0), .S(
        rst), .Z(Red_sel_Key[0]) );
  MUX2_X1 Red_selectsMUX_MUXInst_1_U1 ( .A(Red_selectsReg[1]), .B(1'b0), .S(
        rst), .Z(Red_sel_Key[1]) );
  MUX2_X1 Red_selectsMUX_MUXInst_2_U1 ( .A(Red_selectsReg[2]), .B(1'b0), .S(
        rst), .Z(Red_sel_Key[2]) );
  MUX2_X1 Red_selectsMUX_MUXInst_3_U1 ( .A(Red_selectsReg[3]), .B(1'b0), .S(
        rst), .Z(Red_sel_Tweak[0]) );
  MUX2_X1 Red_selectsMUX_MUXInst_4_U1 ( .A(Red_selectsReg[4]), .B(1'b0), .S(
        rst), .Z(Red_sel_Tweak[1]) );
  MUX2_X1 Red_selectsMUX_MUXInst_5_U1 ( .A(Red_selectsReg[5]), .B(1'b0), .S(
        rst), .Z(Red_sel_Tweak[2]) );
  INV_X1 Red_selectsUpdateInst_Red_selectsUpdateBitInst_0_U2 ( .A(selects[0]), 
        .ZN(Red_selectsNext[0]) );
  INV_X1 Red_selectsUpdateInst_Red_selectsUpdateBitInst_1_U2 ( .A(selects[0]), 
        .ZN(Red_selectsNext[1]) );
  XOR2_X1 Red_selectsUpdateInst_Red_selectsUpdateBitInst_3_U2 ( .A(selects[0]), 
        .B(selects[1]), .Z(Red_selectsNext[3]) );
  XOR2_X1 Red_selectsUpdateInst_Red_selectsUpdateBitInst_4_U2 ( .A(selects[0]), 
        .B(selects[1]), .Z(Red_selectsNext[4]) );
  DFF_X1 Red_selectsRegInst_s_current_state_reg_0_ ( .D(Red_selectsNext[0]), 
        .CK(clk), .Q(Red_selectsReg[0]), .QN() );
  DFF_X1 Red_selectsRegInst_s_current_state_reg_1_ ( .D(Red_selectsNext[1]), 
        .CK(clk), .Q(Red_selectsReg[1]), .QN() );
  DFF_X1 Red_selectsRegInst_s_current_state_reg_2_ ( .D(1'b0), .CK(clk), .Q(
        Red_selectsReg[2]), .QN() );
  DFF_X1 Red_selectsRegInst_s_current_state_reg_3_ ( .D(Red_selectsNext[3]), 
        .CK(clk), .Q(Red_selectsReg[3]), .QN() );
  DFF_X1 Red_selectsRegInst_s_current_state_reg_4_ ( .D(Red_selectsNext[4]), 
        .CK(clk), .Q(Red_selectsReg[4]), .QN() );
  DFF_X1 Red_selectsRegInst_s_current_state_reg_5_ ( .D(1'b0), .CK(clk), .Q(
        Red_selectsReg[5]), .QN() );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_0_LFInst_0_n1), .B(AddRoundKeyOutput[2]), .ZN(
        Red_SignaltoCheck[0]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U1 ( .A(AddRoundKeyOutput[0]), 
        .B(AddRoundKeyOutput[1]), .ZN(Red_ToCheckInst_LFInst_0_LFInst_0_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_0_LFInst_1_n1), .B(AddRoundKeyOutput[3]), .ZN(
        Red_SignaltoCheck[1]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_1_U1 ( .A(AddRoundKeyOutput[0]), 
        .B(AddRoundKeyOutput[1]), .ZN(Red_ToCheckInst_LFInst_0_LFInst_1_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_0_LFInst_2_n1), .B(AddRoundKeyOutput[3]), .ZN(
        Red_SignaltoCheck[2]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_2_U1 ( .A(AddRoundKeyOutput[1]), 
        .B(AddRoundKeyOutput[2]), .ZN(Red_ToCheckInst_LFInst_0_LFInst_2_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_1_LFInst_0_n1), .B(AddRoundKeyOutput[6]), .ZN(
        Red_SignaltoCheck[3]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U1 ( .A(AddRoundKeyOutput[4]), 
        .B(AddRoundKeyOutput[5]), .ZN(Red_ToCheckInst_LFInst_1_LFInst_0_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_1_LFInst_1_n1), .B(AddRoundKeyOutput[7]), .ZN(
        Red_SignaltoCheck[4]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_1_U1 ( .A(AddRoundKeyOutput[4]), 
        .B(AddRoundKeyOutput[5]), .ZN(Red_ToCheckInst_LFInst_1_LFInst_1_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_1_LFInst_2_n1), .B(AddRoundKeyOutput[7]), .ZN(
        Red_SignaltoCheck[5]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_2_U1 ( .A(AddRoundKeyOutput[5]), 
        .B(AddRoundKeyOutput[6]), .ZN(Red_ToCheckInst_LFInst_1_LFInst_2_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_2_LFInst_0_n1), .B(AddRoundKeyOutput[10]), .ZN(
        Red_SignaltoCheck[6]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U1 ( .A(AddRoundKeyOutput[8]), 
        .B(AddRoundKeyOutput[9]), .ZN(Red_ToCheckInst_LFInst_2_LFInst_0_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_2_LFInst_1_n1), .B(AddRoundKeyOutput[11]), .ZN(
        Red_SignaltoCheck[7]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_1_U1 ( .A(AddRoundKeyOutput[8]), 
        .B(AddRoundKeyOutput[9]), .ZN(Red_ToCheckInst_LFInst_2_LFInst_1_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_2_LFInst_2_n1), .B(AddRoundKeyOutput[11]), .ZN(
        Red_SignaltoCheck[8]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_2_U1 ( .A(AddRoundKeyOutput[9]), 
        .B(AddRoundKeyOutput[10]), .ZN(Red_ToCheckInst_LFInst_2_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_3_LFInst_0_n1), .B(AddRoundKeyOutput[14]), .ZN(
        Red_SignaltoCheck[9]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U1 ( .A(AddRoundKeyOutput[12]), 
        .B(AddRoundKeyOutput[13]), .ZN(Red_ToCheckInst_LFInst_3_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_3_LFInst_1_n1), .B(AddRoundKeyOutput[15]), .ZN(
        Red_SignaltoCheck[10]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_1_U1 ( .A(AddRoundKeyOutput[12]), 
        .B(AddRoundKeyOutput[13]), .ZN(Red_ToCheckInst_LFInst_3_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_3_LFInst_2_n1), .B(AddRoundKeyOutput[15]), .ZN(
        Red_SignaltoCheck[11]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_2_U1 ( .A(AddRoundKeyOutput[13]), 
        .B(AddRoundKeyOutput[14]), .ZN(Red_ToCheckInst_LFInst_3_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_4_LFInst_0_n1), .B(AddRoundKeyOutput[18]), .ZN(
        Red_SignaltoCheck[12]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U1 ( .A(AddRoundKeyOutput[16]), 
        .B(AddRoundKeyOutput[17]), .ZN(Red_ToCheckInst_LFInst_4_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_4_LFInst_1_n1), .B(AddRoundKeyOutput[19]), .ZN(
        Red_SignaltoCheck[13]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_1_U1 ( .A(AddRoundKeyOutput[16]), 
        .B(AddRoundKeyOutput[17]), .ZN(Red_ToCheckInst_LFInst_4_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_4_LFInst_2_n1), .B(AddRoundKeyOutput[19]), .ZN(
        Red_SignaltoCheck[14]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_2_U1 ( .A(AddRoundKeyOutput[17]), 
        .B(AddRoundKeyOutput[18]), .ZN(Red_ToCheckInst_LFInst_4_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_5_LFInst_0_n1), .B(AddRoundKeyOutput[22]), .ZN(
        Red_SignaltoCheck[15]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U1 ( .A(AddRoundKeyOutput[20]), 
        .B(AddRoundKeyOutput[21]), .ZN(Red_ToCheckInst_LFInst_5_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_5_LFInst_1_n1), .B(AddRoundKeyOutput[23]), .ZN(
        Red_SignaltoCheck[16]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_1_U1 ( .A(AddRoundKeyOutput[20]), 
        .B(AddRoundKeyOutput[21]), .ZN(Red_ToCheckInst_LFInst_5_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_5_LFInst_2_n1), .B(AddRoundKeyOutput[23]), .ZN(
        Red_SignaltoCheck[17]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_2_U1 ( .A(AddRoundKeyOutput[21]), 
        .B(AddRoundKeyOutput[22]), .ZN(Red_ToCheckInst_LFInst_5_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_6_LFInst_0_n1), .B(AddRoundKeyOutput[26]), .ZN(
        Red_SignaltoCheck[18]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U1 ( .A(AddRoundKeyOutput[24]), 
        .B(AddRoundKeyOutput[25]), .ZN(Red_ToCheckInst_LFInst_6_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_6_LFInst_1_n1), .B(AddRoundKeyOutput[27]), .ZN(
        Red_SignaltoCheck[19]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_1_U1 ( .A(AddRoundKeyOutput[24]), 
        .B(AddRoundKeyOutput[25]), .ZN(Red_ToCheckInst_LFInst_6_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_6_LFInst_2_n1), .B(AddRoundKeyOutput[27]), .ZN(
        Red_SignaltoCheck[20]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_2_U1 ( .A(AddRoundKeyOutput[25]), 
        .B(AddRoundKeyOutput[26]), .ZN(Red_ToCheckInst_LFInst_6_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_7_LFInst_0_n1), .B(AddRoundKeyOutput[30]), .ZN(
        Red_SignaltoCheck[21]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U1 ( .A(AddRoundKeyOutput[28]), 
        .B(AddRoundKeyOutput[29]), .ZN(Red_ToCheckInst_LFInst_7_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_7_LFInst_1_n1), .B(AddRoundKeyOutput[31]), .ZN(
        Red_SignaltoCheck[22]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_1_U1 ( .A(AddRoundKeyOutput[28]), 
        .B(AddRoundKeyOutput[29]), .ZN(Red_ToCheckInst_LFInst_7_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_7_LFInst_2_n1), .B(AddRoundKeyOutput[31]), .ZN(
        Red_SignaltoCheck[23]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_2_U1 ( .A(AddRoundKeyOutput[29]), 
        .B(AddRoundKeyOutput[30]), .ZN(Red_ToCheckInst_LFInst_7_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_8_LFInst_0_n1), .B(AddRoundKeyOutput[34]), .ZN(
        Red_SignaltoCheck[24]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U1 ( .A(AddRoundKeyOutput[32]), 
        .B(AddRoundKeyOutput[33]), .ZN(Red_ToCheckInst_LFInst_8_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_8_LFInst_1_n1), .B(AddRoundKeyOutput[35]), .ZN(
        Red_SignaltoCheck[25]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_1_U1 ( .A(AddRoundKeyOutput[32]), 
        .B(AddRoundKeyOutput[33]), .ZN(Red_ToCheckInst_LFInst_8_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_8_LFInst_2_n1), .B(AddRoundKeyOutput[35]), .ZN(
        Red_SignaltoCheck[26]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_2_U1 ( .A(AddRoundKeyOutput[33]), 
        .B(AddRoundKeyOutput[34]), .ZN(Red_ToCheckInst_LFInst_8_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_9_LFInst_0_n1), .B(AddRoundKeyOutput[38]), .ZN(
        Red_SignaltoCheck[27]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U1 ( .A(AddRoundKeyOutput[36]), 
        .B(AddRoundKeyOutput[37]), .ZN(Red_ToCheckInst_LFInst_9_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_9_LFInst_1_n1), .B(AddRoundKeyOutput[39]), .ZN(
        Red_SignaltoCheck[28]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_1_U1 ( .A(AddRoundKeyOutput[36]), 
        .B(AddRoundKeyOutput[37]), .ZN(Red_ToCheckInst_LFInst_9_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_9_LFInst_2_n1), .B(AddRoundKeyOutput[39]), .ZN(
        Red_SignaltoCheck[29]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_2_U1 ( .A(AddRoundKeyOutput[37]), 
        .B(AddRoundKeyOutput[38]), .ZN(Red_ToCheckInst_LFInst_9_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_10_LFInst_0_n1), .B(AddRoundKeyOutput[42]), 
        .ZN(Red_SignaltoCheck[30]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U1 ( .A(AddRoundKeyOutput[40]), 
        .B(AddRoundKeyOutput[41]), .ZN(Red_ToCheckInst_LFInst_10_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_10_LFInst_1_n1), .B(AddRoundKeyOutput[43]), 
        .ZN(Red_SignaltoCheck[31]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_1_U1 ( .A(AddRoundKeyOutput[40]), 
        .B(AddRoundKeyOutput[41]), .ZN(Red_ToCheckInst_LFInst_10_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_10_LFInst_2_n1), .B(AddRoundKeyOutput[43]), 
        .ZN(Red_SignaltoCheck[32]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_2_U1 ( .A(AddRoundKeyOutput[41]), 
        .B(AddRoundKeyOutput[42]), .ZN(Red_ToCheckInst_LFInst_10_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_11_LFInst_0_n1), .B(AddRoundKeyOutput[46]), 
        .ZN(Red_SignaltoCheck[33]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U1 ( .A(AddRoundKeyOutput[44]), 
        .B(AddRoundKeyOutput[45]), .ZN(Red_ToCheckInst_LFInst_11_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_11_LFInst_1_n1), .B(AddRoundKeyOutput[47]), 
        .ZN(Red_SignaltoCheck[34]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_1_U1 ( .A(AddRoundKeyOutput[44]), 
        .B(AddRoundKeyOutput[45]), .ZN(Red_ToCheckInst_LFInst_11_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_11_LFInst_2_n1), .B(AddRoundKeyOutput[47]), 
        .ZN(Red_SignaltoCheck[35]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_2_U1 ( .A(AddRoundKeyOutput[45]), 
        .B(AddRoundKeyOutput[46]), .ZN(Red_ToCheckInst_LFInst_11_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_12_LFInst_0_n1), .B(AddRoundKeyOutput[50]), 
        .ZN(Red_SignaltoCheck[36]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U1 ( .A(AddRoundKeyOutput[48]), 
        .B(AddRoundKeyOutput[49]), .ZN(Red_ToCheckInst_LFInst_12_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_12_LFInst_1_n1), .B(AddRoundKeyOutput[51]), 
        .ZN(Red_SignaltoCheck[37]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_1_U1 ( .A(AddRoundKeyOutput[48]), 
        .B(AddRoundKeyOutput[49]), .ZN(Red_ToCheckInst_LFInst_12_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_12_LFInst_2_n1), .B(AddRoundKeyOutput[51]), 
        .ZN(Red_SignaltoCheck[38]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_2_U1 ( .A(AddRoundKeyOutput[49]), 
        .B(AddRoundKeyOutput[50]), .ZN(Red_ToCheckInst_LFInst_12_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_13_LFInst_0_n1), .B(AddRoundKeyOutput[54]), 
        .ZN(Red_SignaltoCheck[39]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U1 ( .A(AddRoundKeyOutput[52]), 
        .B(AddRoundKeyOutput[53]), .ZN(Red_ToCheckInst_LFInst_13_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_13_LFInst_1_n1), .B(AddRoundKeyOutput[55]), 
        .ZN(Red_SignaltoCheck[40]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_1_U1 ( .A(AddRoundKeyOutput[52]), 
        .B(AddRoundKeyOutput[53]), .ZN(Red_ToCheckInst_LFInst_13_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_13_LFInst_2_n1), .B(AddRoundKeyOutput[55]), 
        .ZN(Red_SignaltoCheck[41]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_2_U1 ( .A(AddRoundKeyOutput[53]), 
        .B(AddRoundKeyOutput[54]), .ZN(Red_ToCheckInst_LFInst_13_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_14_LFInst_0_n1), .B(AddRoundKeyOutput[58]), 
        .ZN(Red_SignaltoCheck[42]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U1 ( .A(AddRoundKeyOutput[56]), 
        .B(AddRoundKeyOutput[57]), .ZN(Red_ToCheckInst_LFInst_14_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_14_LFInst_1_n1), .B(AddRoundKeyOutput[59]), 
        .ZN(Red_SignaltoCheck[43]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_1_U1 ( .A(AddRoundKeyOutput[56]), 
        .B(AddRoundKeyOutput[57]), .ZN(Red_ToCheckInst_LFInst_14_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_14_LFInst_2_n1), .B(AddRoundKeyOutput[59]), 
        .ZN(Red_SignaltoCheck[44]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_2_U1 ( .A(AddRoundKeyOutput[57]), 
        .B(AddRoundKeyOutput[58]), .ZN(Red_ToCheckInst_LFInst_14_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_15_LFInst_0_n1), .B(AddRoundKeyOutput[62]), 
        .ZN(Red_SignaltoCheck[45]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U1 ( .A(AddRoundKeyOutput[60]), 
        .B(AddRoundKeyOutput[61]), .ZN(Red_ToCheckInst_LFInst_15_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_15_LFInst_1_n1), .B(AddRoundKeyOutput[63]), 
        .ZN(Red_SignaltoCheck[46]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_1_U1 ( .A(AddRoundKeyOutput[60]), 
        .B(AddRoundKeyOutput[61]), .ZN(Red_ToCheckInst_LFInst_15_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_15_LFInst_2_n1), .B(AddRoundKeyOutput[63]), 
        .ZN(Red_SignaltoCheck[47]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_2_U1 ( .A(AddRoundKeyOutput[61]), 
        .B(AddRoundKeyOutput[62]), .ZN(Red_ToCheckInst_LFInst_15_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_16_LFInst_0_n1), .B(FSMUpdate[2]), .ZN(
        Red_SignaltoCheck[48]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U1 ( .A(FSMUpdate[0]), .B(
        FSMUpdate[1]), .ZN(Red_ToCheckInst_LFInst_16_LFInst_0_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_16_LFInst_1_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[49]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_1_U1 ( .A(FSMUpdate[0]), .B(
        FSMUpdate[1]), .ZN(Red_ToCheckInst_LFInst_16_LFInst_1_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_16_LFInst_2_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[50]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_2_U1 ( .A(FSMUpdate[1]), .B(
        FSMUpdate[2]), .ZN(Red_ToCheckInst_LFInst_16_LFInst_2_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_17_LFInst_0_n1), .B(FSMUpdate[5]), .ZN(
        Red_SignaltoCheck[51]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U1 ( .A(FSMUpdate[3]), .B(
        FSMUpdate[4]), .ZN(Red_ToCheckInst_LFInst_17_LFInst_0_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_17_LFInst_1_n1), .B(FSMUpdate[6]), .ZN(
        Red_SignaltoCheck[52]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_1_U1 ( .A(FSMUpdate[3]), .B(
        FSMUpdate[4]), .ZN(Red_ToCheckInst_LFInst_17_LFInst_1_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_17_LFInst_2_n1), .B(FSMUpdate[6]), .ZN(
        Red_SignaltoCheck[53]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_2_U1 ( .A(FSMUpdate[4]), .B(
        FSMUpdate[5]), .ZN(Red_ToCheckInst_LFInst_17_LFInst_2_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_18_LFInst_0_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[54]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U1 ( .A(selectsNext[0]), .B(1'b0), .ZN(Red_ToCheckInst_LFInst_18_LFInst_0_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_18_LFInst_1_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[55]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_1_U1 ( .A(selectsNext[0]), .B(1'b0), .ZN(Red_ToCheckInst_LFInst_18_LFInst_1_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_18_LFInst_2_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[56]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_2_U1 ( .A(1'b0), .B(1'b0), .ZN(
        Red_ToCheckInst_LFInst_18_LFInst_2_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_19_LFInst_0_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[57]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U1 ( .A(selectsNext[1]), .B(1'b0), .ZN(Red_ToCheckInst_LFInst_19_LFInst_0_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_19_LFInst_1_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[58]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_1_U1 ( .A(selectsNext[1]), .B(1'b0), .ZN(Red_ToCheckInst_LFInst_19_LFInst_1_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_19_LFInst_2_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[59]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_2_U1 ( .A(1'b0), .B(1'b0), .ZN(
        Red_ToCheckInst_LFInst_19_LFInst_2_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_20_LFInst_0_n1), .B(PermutationOutput[62]), 
        .ZN(Red_SignaltoCheck[60]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U1 ( .A(PermutationOutput[60]), 
        .B(PermutationOutput[61]), .ZN(Red_ToCheckInst_LFInst_20_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_20_LFInst_1_n1), .B(PermutationOutput[63]), 
        .ZN(Red_SignaltoCheck[61]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_1_U1 ( .A(PermutationOutput[60]), 
        .B(PermutationOutput[61]), .ZN(Red_ToCheckInst_LFInst_20_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_20_LFInst_2_n1), .B(PermutationOutput[63]), 
        .ZN(Red_SignaltoCheck[62]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_2_U1 ( .A(PermutationOutput[61]), 
        .B(PermutationOutput[62]), .ZN(Red_ToCheckInst_LFInst_20_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_21_LFInst_0_n1), .B(PermutationOutput[50]), 
        .ZN(Red_SignaltoCheck[63]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U1 ( .A(PermutationOutput[48]), 
        .B(PermutationOutput[49]), .ZN(Red_ToCheckInst_LFInst_21_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_21_LFInst_1_n1), .B(PermutationOutput[51]), 
        .ZN(Red_SignaltoCheck[64]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_1_U1 ( .A(PermutationOutput[48]), 
        .B(PermutationOutput[49]), .ZN(Red_ToCheckInst_LFInst_21_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_21_LFInst_2_n1), .B(PermutationOutput[51]), 
        .ZN(Red_SignaltoCheck[65]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_2_U1 ( .A(PermutationOutput[49]), 
        .B(PermutationOutput[50]), .ZN(Red_ToCheckInst_LFInst_21_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_22_LFInst_0_n1), .B(PermutationOutput[54]), 
        .ZN(Red_SignaltoCheck[66]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U1 ( .A(PermutationOutput[52]), 
        .B(PermutationOutput[53]), .ZN(Red_ToCheckInst_LFInst_22_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_22_LFInst_1_n1), .B(PermutationOutput[55]), 
        .ZN(Red_SignaltoCheck[67]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_1_U1 ( .A(PermutationOutput[52]), 
        .B(PermutationOutput[53]), .ZN(Red_ToCheckInst_LFInst_22_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_22_LFInst_2_n1), .B(PermutationOutput[55]), 
        .ZN(Red_SignaltoCheck[68]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_2_U1 ( .A(PermutationOutput[53]), 
        .B(PermutationOutput[54]), .ZN(Red_ToCheckInst_LFInst_22_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_23_LFInst_0_n1), .B(PermutationOutput[58]), 
        .ZN(Red_SignaltoCheck[69]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U1 ( .A(PermutationOutput[56]), 
        .B(PermutationOutput[57]), .ZN(Red_ToCheckInst_LFInst_23_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_23_LFInst_1_n1), .B(PermutationOutput[59]), 
        .ZN(Red_SignaltoCheck[70]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_1_U1 ( .A(PermutationOutput[56]), 
        .B(PermutationOutput[57]), .ZN(Red_ToCheckInst_LFInst_23_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_23_LFInst_2_n1), .B(PermutationOutput[59]), 
        .ZN(Red_SignaltoCheck[71]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_2_U1 ( .A(PermutationOutput[57]), 
        .B(PermutationOutput[58]), .ZN(Red_ToCheckInst_LFInst_23_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_24_LFInst_0_n1), .B(PermutationOutput[34]), 
        .ZN(Red_SignaltoCheck[72]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U1 ( .A(PermutationOutput[32]), 
        .B(PermutationOutput[33]), .ZN(Red_ToCheckInst_LFInst_24_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_24_LFInst_1_n1), .B(PermutationOutput[35]), 
        .ZN(Red_SignaltoCheck[73]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_1_U1 ( .A(PermutationOutput[32]), 
        .B(PermutationOutput[33]), .ZN(Red_ToCheckInst_LFInst_24_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_24_LFInst_2_n1), .B(PermutationOutput[35]), 
        .ZN(Red_SignaltoCheck[74]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_2_U1 ( .A(PermutationOutput[33]), 
        .B(PermutationOutput[34]), .ZN(Red_ToCheckInst_LFInst_24_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_25_LFInst_0_n1), .B(PermutationOutput[46]), 
        .ZN(Red_SignaltoCheck[75]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U1 ( .A(PermutationOutput[44]), 
        .B(PermutationOutput[45]), .ZN(Red_ToCheckInst_LFInst_25_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_25_LFInst_1_n1), .B(PermutationOutput[47]), 
        .ZN(Red_SignaltoCheck[76]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_1_U1 ( .A(PermutationOutput[44]), 
        .B(PermutationOutput[45]), .ZN(Red_ToCheckInst_LFInst_25_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_25_LFInst_2_n1), .B(PermutationOutput[47]), 
        .ZN(Red_SignaltoCheck[77]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_2_U1 ( .A(PermutationOutput[45]), 
        .B(PermutationOutput[46]), .ZN(Red_ToCheckInst_LFInst_25_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_26_LFInst_0_n1), .B(PermutationOutput[42]), 
        .ZN(Red_SignaltoCheck[78]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U1 ( .A(PermutationOutput[40]), 
        .B(PermutationOutput[41]), .ZN(Red_ToCheckInst_LFInst_26_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_26_LFInst_1_n1), .B(PermutationOutput[43]), 
        .ZN(Red_SignaltoCheck[79]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_1_U1 ( .A(PermutationOutput[40]), 
        .B(PermutationOutput[41]), .ZN(Red_ToCheckInst_LFInst_26_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_26_LFInst_2_n1), .B(PermutationOutput[43]), 
        .ZN(Red_SignaltoCheck[80]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_2_U1 ( .A(PermutationOutput[41]), 
        .B(PermutationOutput[42]), .ZN(Red_ToCheckInst_LFInst_26_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_27_LFInst_0_n1), .B(PermutationOutput[38]), 
        .ZN(Red_SignaltoCheck[81]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U1 ( .A(PermutationOutput[36]), 
        .B(PermutationOutput[37]), .ZN(Red_ToCheckInst_LFInst_27_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_27_LFInst_1_n1), .B(PermutationOutput[39]), 
        .ZN(Red_SignaltoCheck[82]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_1_U1 ( .A(PermutationOutput[36]), 
        .B(PermutationOutput[37]), .ZN(Red_ToCheckInst_LFInst_27_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_27_LFInst_2_n1), .B(PermutationOutput[39]), 
        .ZN(Red_SignaltoCheck[83]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_2_U1 ( .A(PermutationOutput[37]), 
        .B(PermutationOutput[38]), .ZN(Red_ToCheckInst_LFInst_27_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_28_LFInst_0_n1), .B(PermutationOutput[18]), 
        .ZN(Red_SignaltoCheck[84]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U1 ( .A(PermutationOutput[16]), 
        .B(PermutationOutput[17]), .ZN(Red_ToCheckInst_LFInst_28_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_28_LFInst_1_n1), .B(PermutationOutput[19]), 
        .ZN(Red_SignaltoCheck[85]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_1_U1 ( .A(PermutationOutput[16]), 
        .B(PermutationOutput[17]), .ZN(Red_ToCheckInst_LFInst_28_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_28_LFInst_2_n1), .B(PermutationOutput[19]), 
        .ZN(Red_SignaltoCheck[86]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_2_U1 ( .A(PermutationOutput[17]), 
        .B(PermutationOutput[18]), .ZN(Red_ToCheckInst_LFInst_28_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_29_LFInst_0_n1), .B(PermutationOutput[30]), 
        .ZN(Red_SignaltoCheck[87]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U1 ( .A(PermutationOutput[28]), 
        .B(PermutationOutput[29]), .ZN(Red_ToCheckInst_LFInst_29_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_29_LFInst_1_n1), .B(PermutationOutput[31]), 
        .ZN(Red_SignaltoCheck[88]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_1_U1 ( .A(PermutationOutput[28]), 
        .B(PermutationOutput[29]), .ZN(Red_ToCheckInst_LFInst_29_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_29_LFInst_2_n1), .B(PermutationOutput[31]), 
        .ZN(Red_SignaltoCheck[89]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_2_U1 ( .A(PermutationOutput[29]), 
        .B(PermutationOutput[30]), .ZN(Red_ToCheckInst_LFInst_29_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_30_LFInst_0_n1), .B(PermutationOutput[26]), 
        .ZN(Red_SignaltoCheck[90]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U1 ( .A(PermutationOutput[24]), 
        .B(PermutationOutput[25]), .ZN(Red_ToCheckInst_LFInst_30_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_30_LFInst_1_n1), .B(PermutationOutput[27]), 
        .ZN(Red_SignaltoCheck[91]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_1_U1 ( .A(PermutationOutput[24]), 
        .B(PermutationOutput[25]), .ZN(Red_ToCheckInst_LFInst_30_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_30_LFInst_2_n1), .B(PermutationOutput[27]), 
        .ZN(Red_SignaltoCheck[92]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_2_U1 ( .A(PermutationOutput[25]), 
        .B(PermutationOutput[26]), .ZN(Red_ToCheckInst_LFInst_30_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_31_LFInst_0_n1), .B(PermutationOutput[22]), 
        .ZN(Red_SignaltoCheck[93]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U1 ( .A(PermutationOutput[20]), 
        .B(PermutationOutput[21]), .ZN(Red_ToCheckInst_LFInst_31_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_31_LFInst_1_n1), .B(PermutationOutput[23]), 
        .ZN(Red_SignaltoCheck[94]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_1_U1 ( .A(PermutationOutput[20]), 
        .B(PermutationOutput[21]), .ZN(Red_ToCheckInst_LFInst_31_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_31_LFInst_2_n1), .B(PermutationOutput[23]), 
        .ZN(Red_SignaltoCheck[95]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_2_U1 ( .A(PermutationOutput[21]), 
        .B(PermutationOutput[22]), .ZN(Red_ToCheckInst_LFInst_31_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_32_LFInst_0_n1), .B(PermutationOutput[6]), .ZN(
        Red_SignaltoCheck[96]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U1 ( .A(PermutationOutput[4]), 
        .B(PermutationOutput[5]), .ZN(Red_ToCheckInst_LFInst_32_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_32_LFInst_1_n1), .B(PermutationOutput[7]), .ZN(
        Red_SignaltoCheck[97]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_1_U1 ( .A(PermutationOutput[4]), 
        .B(PermutationOutput[5]), .ZN(Red_ToCheckInst_LFInst_32_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_32_LFInst_2_n1), .B(PermutationOutput[7]), .ZN(
        Red_SignaltoCheck[98]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_2_U1 ( .A(PermutationOutput[5]), 
        .B(PermutationOutput[6]), .ZN(Red_ToCheckInst_LFInst_32_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_33_LFInst_0_n1), .B(PermutationOutput[10]), 
        .ZN(Red_SignaltoCheck[99]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U1 ( .A(PermutationOutput[8]), 
        .B(PermutationOutput[9]), .ZN(Red_ToCheckInst_LFInst_33_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_33_LFInst_1_n1), .B(PermutationOutput[11]), 
        .ZN(Red_SignaltoCheck[100]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_1_U1 ( .A(PermutationOutput[8]), 
        .B(PermutationOutput[9]), .ZN(Red_ToCheckInst_LFInst_33_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_33_LFInst_2_n1), .B(PermutationOutput[11]), 
        .ZN(Red_SignaltoCheck[101]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_2_U1 ( .A(PermutationOutput[9]), 
        .B(PermutationOutput[10]), .ZN(Red_ToCheckInst_LFInst_33_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_34_LFInst_0_n1), .B(PermutationOutput[14]), 
        .ZN(Red_SignaltoCheck[102]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U1 ( .A(PermutationOutput[12]), 
        .B(PermutationOutput[13]), .ZN(Red_ToCheckInst_LFInst_34_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_34_LFInst_1_n1), .B(PermutationOutput[15]), 
        .ZN(Red_SignaltoCheck[103]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_1_U1 ( .A(PermutationOutput[12]), 
        .B(PermutationOutput[13]), .ZN(Red_ToCheckInst_LFInst_34_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_34_LFInst_2_n1), .B(PermutationOutput[15]), 
        .ZN(Red_SignaltoCheck[104]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_2_U1 ( .A(PermutationOutput[13]), 
        .B(PermutationOutput[14]), .ZN(Red_ToCheckInst_LFInst_34_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_35_LFInst_0_n1), .B(PermutationOutput[2]), .ZN(
        Red_SignaltoCheck[105]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U1 ( .A(PermutationOutput[0]), 
        .B(PermutationOutput[1]), .ZN(Red_ToCheckInst_LFInst_35_LFInst_0_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_35_LFInst_1_n1), .B(PermutationOutput[3]), .ZN(
        Red_SignaltoCheck[106]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_1_U1 ( .A(PermutationOutput[0]), 
        .B(PermutationOutput[1]), .ZN(Red_ToCheckInst_LFInst_35_LFInst_1_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_35_LFInst_2_n1), .B(PermutationOutput[3]), .ZN(
        Red_SignaltoCheck[107]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_2_U1 ( .A(PermutationOutput[1]), 
        .B(PermutationOutput[2]), .ZN(Red_ToCheckInst_LFInst_35_LFInst_2_n1)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_36_LFInst_0_n1), .B(FSMUpdate[1]), .ZN(
        Red_SignaltoCheck[108]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U1 ( .A(RoundConstant_0), .B(
        FSMUpdate[0]), .ZN(Red_ToCheckInst_LFInst_36_LFInst_0_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_36_LFInst_1_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[109]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_1_U1 ( .A(RoundConstant_0), .B(
        FSMUpdate[0]), .ZN(Red_ToCheckInst_LFInst_36_LFInst_1_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_36_LFInst_2_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[110]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_2_U1 ( .A(FSMUpdate[0]), .B(
        FSMUpdate[1]), .ZN(Red_ToCheckInst_LFInst_36_LFInst_2_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_37_LFInst_0_n1), .B(FSMUpdate[4]), .ZN(
        Red_SignaltoCheck[111]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U1 ( .A(RoundConstant_4_), .B(
        FSMUpdate[3]), .ZN(Red_ToCheckInst_LFInst_37_LFInst_0_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_37_LFInst_1_n1), .B(FSMUpdate[5]), .ZN(
        Red_SignaltoCheck[112]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_1_U1 ( .A(RoundConstant_4_), .B(
        FSMUpdate[3]), .ZN(Red_ToCheckInst_LFInst_37_LFInst_1_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_37_LFInst_2_n1), .B(FSMUpdate[5]), .ZN(
        Red_SignaltoCheck[113]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_2_U1 ( .A(FSMUpdate[3]), .B(
        FSMUpdate[4]), .ZN(Red_ToCheckInst_LFInst_37_LFInst_2_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_38_LFInst_0_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[114]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U1 ( .A(selects[1]), .B(1'b0), 
        .ZN(Red_ToCheckInst_LFInst_38_LFInst_0_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_38_LFInst_1_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[115]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_1_U1 ( .A(selects[1]), .B(1'b0), 
        .ZN(Red_ToCheckInst_LFInst_38_LFInst_1_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_38_LFInst_2_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[116]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_2_U1 ( .A(1'b0), .B(1'b0), .ZN(
        Red_ToCheckInst_LFInst_38_LFInst_2_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_39_LFInst_0_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[117]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U1 ( .A(selects[0]), .B(1'b0), 
        .ZN(Red_ToCheckInst_LFInst_39_LFInst_0_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_39_LFInst_1_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[118]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_1_U1 ( .A(selects[0]), .B(1'b0), 
        .ZN(Red_ToCheckInst_LFInst_39_LFInst_1_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_39_LFInst_2_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[119]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_2_U1 ( .A(1'b0), .B(1'b0), .ZN(
        Red_ToCheckInst_LFInst_39_LFInst_2_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U2 ( .A(
        Red_ToCheckInst_LFInst_40_LFInst_0_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[120]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U1 ( .A(done), .B(1'b0), .ZN(
        Red_ToCheckInst_LFInst_40_LFInst_0_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_1_U2 ( .A(
        Red_ToCheckInst_LFInst_40_LFInst_1_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[121]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_1_U1 ( .A(done), .B(1'b0), .ZN(
        Red_ToCheckInst_LFInst_40_LFInst_1_n1) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_2_U2 ( .A(
        Red_ToCheckInst_LFInst_40_LFInst_2_n1), .B(1'b0), .ZN(
        Red_SignaltoCheck[122]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_2_U1 ( .A(1'b0), .B(1'b0), .ZN(
        Red_ToCheckInst_LFInst_40_LFInst_2_n1) );
  NAND4_X1 Check1_CheckInst_0_U55 ( .A1(Check1_CheckInst_0_n52), .A2(
        Check1_CheckInst_0_n51), .A3(Check1_CheckInst_0_n50), .A4(
        Check1_CheckInst_0_n49), .ZN(Check1_CheckInst_0_n53) );
  XNOR2_X1 Check1_CheckInst_0_U54 ( .A(Red_StateRegOutput[36]), .B(
        Red_SignaltoCheck[96]), .ZN(Check1_CheckInst_0_n49) );
  XNOR2_X1 Check1_CheckInst_0_U53 ( .A(Red_done[0]), .B(Red_SignaltoCheck[120]), .ZN(Check1_CheckInst_0_n50) );
  NOR4_X1 Check1_CheckInst_0_U52 ( .A1(Check1_CheckInst_0_n48), .A2(
        Check1_CheckInst_0_n47), .A3(Check1_CheckInst_0_n46), .A4(
        Check1_CheckInst_0_n45), .ZN(Check1_CheckInst_0_n51) );
  NAND4_X1 Check1_CheckInst_0_U51 ( .A1(Check1_CheckInst_0_n44), .A2(
        Check1_CheckInst_0_n43), .A3(Check1_CheckInst_0_n42), .A4(
        Check1_CheckInst_0_n41), .ZN(Check1_CheckInst_0_n45) );
  NOR4_X1 Check1_CheckInst_0_U50 ( .A1(Check1_CheckInst_0_n40), .A2(
        Check1_CheckInst_0_n39), .A3(Check1_CheckInst_0_n38), .A4(
        Check1_CheckInst_0_n37), .ZN(Check1_CheckInst_0_n41) );
  XOR2_X1 Check1_CheckInst_0_U49 ( .A(Red_final[42]), .B(Red_SignaltoCheck[42]), .Z(Check1_CheckInst_0_n37) );
  XOR2_X1 Check1_CheckInst_0_U48 ( .A(Red_final[33]), .B(Red_SignaltoCheck[33]), .Z(Check1_CheckInst_0_n38) );
  XOR2_X1 Check1_CheckInst_0_U47 ( .A(Red_final[39]), .B(Red_SignaltoCheck[39]), .Z(Check1_CheckInst_0_n39) );
  XOR2_X1 Check1_CheckInst_0_U46 ( .A(Red_final[36]), .B(Red_SignaltoCheck[36]), .Z(Check1_CheckInst_0_n40) );
  NOR4_X1 Check1_CheckInst_0_U45 ( .A1(Check1_CheckInst_0_n36), .A2(
        Check1_CheckInst_0_n35), .A3(Check1_CheckInst_0_n34), .A4(
        Check1_CheckInst_0_n33), .ZN(Check1_CheckInst_0_n42) );
  XOR2_X1 Check1_CheckInst_0_U44 ( .A(Red_final[30]), .B(Red_SignaltoCheck[30]), .Z(Check1_CheckInst_0_n33) );
  XOR2_X1 Check1_CheckInst_0_U43 ( .A(Red_final[27]), .B(Red_SignaltoCheck[27]), .Z(Check1_CheckInst_0_n34) );
  XOR2_X1 Check1_CheckInst_0_U42 ( .A(Red_final[18]), .B(Red_SignaltoCheck[18]), .Z(Check1_CheckInst_0_n35) );
  XOR2_X1 Check1_CheckInst_0_U41 ( .A(Red_final[24]), .B(Red_SignaltoCheck[24]), .Z(Check1_CheckInst_0_n36) );
  NOR4_X1 Check1_CheckInst_0_U40 ( .A1(Check1_CheckInst_0_n32), .A2(
        Check1_CheckInst_0_n31), .A3(Check1_CheckInst_0_n30), .A4(
        Check1_CheckInst_0_n29), .ZN(Check1_CheckInst_0_n43) );
  XOR2_X1 Check1_CheckInst_0_U39 ( .A(Red_final[21]), .B(Red_SignaltoCheck[21]), .Z(Check1_CheckInst_0_n29) );
  XOR2_X1 Check1_CheckInst_0_U38 ( .A(Red_sel_Tweak[0]), .B(
        Red_SignaltoCheck[114]), .Z(Check1_CheckInst_0_n30) );
  XOR2_X1 Check1_CheckInst_0_U37 ( .A(Red_SignaltoCheck[105]), .B(
        Red_StateRegOutput[45]), .Z(Check1_CheckInst_0_n31) );
  XOR2_X1 Check1_CheckInst_0_U36 ( .A(Red_SignaltoCheck[12]), .B(Red_final[12]), .Z(Check1_CheckInst_0_n32) );
  NOR4_X1 Check1_CheckInst_0_U35 ( .A1(Check1_CheckInst_0_n28), .A2(
        Check1_CheckInst_0_n27), .A3(Check1_CheckInst_0_n26), .A4(
        Check1_CheckInst_0_n25), .ZN(Check1_CheckInst_0_n44) );
  XOR2_X1 Check1_CheckInst_0_U34 ( .A(Red_sel_Key[0]), .B(
        Red_SignaltoCheck[117]), .Z(Check1_CheckInst_0_n25) );
  XOR2_X1 Check1_CheckInst_0_U33 ( .A(Red_RoundConstant[3]), .B(
        Red_SignaltoCheck[111]), .Z(Check1_CheckInst_0_n26) );
  XOR2_X1 Check1_CheckInst_0_U32 ( .A(Red_final[0]), .B(Red_SignaltoCheck[0]), 
        .Z(Check1_CheckInst_0_n27) );
  XOR2_X1 Check1_CheckInst_0_U31 ( .A(Red_StateRegOutput[42]), .B(
        Red_SignaltoCheck[102]), .Z(Check1_CheckInst_0_n28) );
  NAND4_X1 Check1_CheckInst_0_U30 ( .A1(Check1_CheckInst_0_n24), .A2(
        Check1_CheckInst_0_n23), .A3(Check1_CheckInst_0_n22), .A4(
        Check1_CheckInst_0_n21), .ZN(Check1_CheckInst_0_n46) );
  XNOR2_X1 Check1_CheckInst_0_U29 ( .A(Red_final[9]), .B(Red_SignaltoCheck[9]), 
        .ZN(Check1_CheckInst_0_n21) );
  XNOR2_X1 Check1_CheckInst_0_U28 ( .A(Red_StateRegOutput[15]), .B(
        Red_SignaltoCheck[75]), .ZN(Check1_CheckInst_0_n22) );
  XNOR2_X1 Check1_CheckInst_0_U27 ( .A(Red_RoundConstant[0]), .B(
        Red_SignaltoCheck[108]), .ZN(Check1_CheckInst_0_n23) );
  NOR4_X1 Check1_CheckInst_0_U26 ( .A1(Check1_CheckInst_0_n20), .A2(
        Check1_CheckInst_0_n19), .A3(Check1_CheckInst_0_n18), .A4(
        Check1_CheckInst_0_n17), .ZN(Check1_CheckInst_0_n24) );
  XOR2_X1 Check1_CheckInst_0_U25 ( .A(Red_final[15]), .B(Red_SignaltoCheck[15]), .Z(Check1_CheckInst_0_n17) );
  XOR2_X1 Check1_CheckInst_0_U24 ( .A(Red_StateRegOutput[18]), .B(
        Red_SignaltoCheck[78]), .Z(Check1_CheckInst_0_n18) );
  XOR2_X1 Check1_CheckInst_0_U23 ( .A(Red_StateRegOutput[12]), .B(
        Red_SignaltoCheck[72]), .Z(Check1_CheckInst_0_n19) );
  XOR2_X1 Check1_CheckInst_0_U22 ( .A(Red_StateRegOutput[27]), .B(
        Red_SignaltoCheck[87]), .Z(Check1_CheckInst_0_n20) );
  XOR2_X1 Check1_CheckInst_0_U21 ( .A(Red_StateRegOutput[3]), .B(
        Red_SignaltoCheck[63]), .Z(Check1_CheckInst_0_n47) );
  XOR2_X1 Check1_CheckInst_0_U20 ( .A(Red_FSMUpdate[0]), .B(
        Red_SignaltoCheck[48]), .Z(Check1_CheckInst_0_n48) );
  NOR3_X1 Check1_CheckInst_0_U19 ( .A1(Check1_CheckInst_0_n16), .A2(
        Check1_CheckInst_0_n15), .A3(Check1_CheckInst_0_n14), .ZN(
        Check1_CheckInst_0_n52) );
  NAND4_X1 Check1_CheckInst_0_U18 ( .A1(Check1_CheckInst_0_n13), .A2(
        Check1_CheckInst_0_n12), .A3(Check1_CheckInst_0_n11), .A4(
        Check1_CheckInst_0_n10), .ZN(Check1_CheckInst_0_n14) );
  XNOR2_X1 Check1_CheckInst_0_U17 ( .A(Red_selectsNext[3]), .B(
        Red_SignaltoCheck[57]), .ZN(Check1_CheckInst_0_n10) );
  XNOR2_X1 Check1_CheckInst_0_U16 ( .A(Red_StateRegOutput[24]), .B(
        Red_SignaltoCheck[84]), .ZN(Check1_CheckInst_0_n11) );
  XNOR2_X1 Check1_CheckInst_0_U15 ( .A(Red_StateRegOutput[9]), .B(
        Red_SignaltoCheck[69]), .ZN(Check1_CheckInst_0_n12) );
  XNOR2_X1 Check1_CheckInst_0_U14 ( .A(Red_StateRegOutput[21]), .B(
        Red_SignaltoCheck[81]), .ZN(Check1_CheckInst_0_n13) );
  XOR2_X1 Check1_CheckInst_0_U13 ( .A(Red_final[3]), .B(Red_SignaltoCheck[3]), 
        .Z(Check1_CheckInst_0_n15) );
  XOR2_X1 Check1_CheckInst_0_U12 ( .A(Red_SignaltoCheck[6]), .B(Red_final[6]), 
        .Z(Check1_CheckInst_0_n16) );
  XNOR2_X1 Check1_CheckInst_0_U11 ( .A(Red_StateRegOutput[0]), .B(
        Red_SignaltoCheck[60]), .ZN(Check1_CheckInst_0_n7) );
  XNOR2_X1 Check1_CheckInst_0_U10 ( .A(Red_SignaltoCheck[66]), .B(
        Red_StateRegOutput[6]), .ZN(Check1_CheckInst_0_n8) );
  NOR4_X1 Check1_CheckInst_0_U9 ( .A1(Check1_CheckInst_0_n6), .A2(
        Check1_CheckInst_0_n5), .A3(Check1_CheckInst_0_n4), .A4(
        Check1_CheckInst_0_n3), .ZN(Check1_CheckInst_0_n9) );
  XOR2_X1 Check1_CheckInst_0_U8 ( .A(Red_StateRegOutput[33]), .B(
        Red_SignaltoCheck[93]), .Z(Check1_CheckInst_0_n3) );
  XOR2_X1 Check1_CheckInst_0_U7 ( .A(Red_StateRegOutput[39]), .B(
        Red_SignaltoCheck[99]), .Z(Check1_CheckInst_0_n4) );
  XOR2_X1 Check1_CheckInst_0_U6 ( .A(Red_selectsNext[0]), .B(
        Red_SignaltoCheck[54]), .Z(Check1_CheckInst_0_n5) );
  XOR2_X1 Check1_CheckInst_0_U5 ( .A(Red_StateRegOutput[30]), .B(
        Red_SignaltoCheck[90]), .Z(Check1_CheckInst_0_n6) );
  XOR2_X1 Check1_CheckInst_0_U4 ( .A(Red_final[45]), .B(Red_SignaltoCheck[45]), 
        .Z(Check1_CheckInst_0_n54) );
  NOR3_X1 Check1_CheckInst_0_U3 ( .A1(Check1_CheckInst_0_n54), .A2(
        Check1_CheckInst_0_n53), .A3(Check1_CheckInst_0_n2), .ZN(Error[0]) );
  NAND4_X1 Check1_CheckInst_0_U2 ( .A1(Check1_CheckInst_0_n9), .A2(
        Check1_CheckInst_0_n7), .A3(Check1_CheckInst_0_n8), .A4(
        Check1_CheckInst_0_n1), .ZN(Check1_CheckInst_0_n2) );
  XNOR2_X1 Check1_CheckInst_0_U1 ( .A(Red_FSMUpdate[3]), .B(
        Red_SignaltoCheck[51]), .ZN(Check1_CheckInst_0_n1) );
  NAND4_X1 Check1_CheckInst_1_U55 ( .A1(Check1_CheckInst_1_n52), .A2(
        Check1_CheckInst_1_n51), .A3(Check1_CheckInst_1_n50), .A4(
        Check1_CheckInst_1_n49), .ZN(Check1_CheckInst_1_n53) );
  XNOR2_X1 Check1_CheckInst_1_U54 ( .A(Red_StateRegOutput[37]), .B(
        Red_SignaltoCheck[97]), .ZN(Check1_CheckInst_1_n49) );
  XNOR2_X1 Check1_CheckInst_1_U53 ( .A(Red_done[1]), .B(Red_SignaltoCheck[121]), .ZN(Check1_CheckInst_1_n50) );
  NOR4_X1 Check1_CheckInst_1_U52 ( .A1(Check1_CheckInst_1_n48), .A2(
        Check1_CheckInst_1_n47), .A3(Check1_CheckInst_1_n46), .A4(
        Check1_CheckInst_1_n45), .ZN(Check1_CheckInst_1_n51) );
  NAND4_X1 Check1_CheckInst_1_U51 ( .A1(Check1_CheckInst_1_n44), .A2(
        Check1_CheckInst_1_n43), .A3(Check1_CheckInst_1_n42), .A4(
        Check1_CheckInst_1_n41), .ZN(Check1_CheckInst_1_n45) );
  NOR4_X1 Check1_CheckInst_1_U50 ( .A1(Check1_CheckInst_1_n40), .A2(
        Check1_CheckInst_1_n39), .A3(Check1_CheckInst_1_n38), .A4(
        Check1_CheckInst_1_n37), .ZN(Check1_CheckInst_1_n41) );
  XOR2_X1 Check1_CheckInst_1_U49 ( .A(Red_final[43]), .B(Red_SignaltoCheck[43]), .Z(Check1_CheckInst_1_n37) );
  XOR2_X1 Check1_CheckInst_1_U48 ( .A(Red_final[34]), .B(Red_SignaltoCheck[34]), .Z(Check1_CheckInst_1_n38) );
  XOR2_X1 Check1_CheckInst_1_U47 ( .A(Red_final[40]), .B(Red_SignaltoCheck[40]), .Z(Check1_CheckInst_1_n39) );
  XOR2_X1 Check1_CheckInst_1_U46 ( .A(Red_final[37]), .B(Red_SignaltoCheck[37]), .Z(Check1_CheckInst_1_n40) );
  NOR4_X1 Check1_CheckInst_1_U45 ( .A1(Check1_CheckInst_1_n36), .A2(
        Check1_CheckInst_1_n35), .A3(Check1_CheckInst_1_n34), .A4(
        Check1_CheckInst_1_n33), .ZN(Check1_CheckInst_1_n42) );
  XOR2_X1 Check1_CheckInst_1_U44 ( .A(Red_final[31]), .B(Red_SignaltoCheck[31]), .Z(Check1_CheckInst_1_n33) );
  XOR2_X1 Check1_CheckInst_1_U43 ( .A(Red_final[28]), .B(Red_SignaltoCheck[28]), .Z(Check1_CheckInst_1_n34) );
  XOR2_X1 Check1_CheckInst_1_U42 ( .A(Red_final[19]), .B(Red_SignaltoCheck[19]), .Z(Check1_CheckInst_1_n35) );
  XOR2_X1 Check1_CheckInst_1_U41 ( .A(Red_final[25]), .B(Red_SignaltoCheck[25]), .Z(Check1_CheckInst_1_n36) );
  NOR4_X1 Check1_CheckInst_1_U40 ( .A1(Check1_CheckInst_1_n32), .A2(
        Check1_CheckInst_1_n31), .A3(Check1_CheckInst_1_n30), .A4(
        Check1_CheckInst_1_n29), .ZN(Check1_CheckInst_1_n43) );
  XOR2_X1 Check1_CheckInst_1_U39 ( .A(Red_final[22]), .B(Red_SignaltoCheck[22]), .Z(Check1_CheckInst_1_n29) );
  XOR2_X1 Check1_CheckInst_1_U38 ( .A(Red_sel_Tweak[1]), .B(
        Red_SignaltoCheck[115]), .Z(Check1_CheckInst_1_n30) );
  XOR2_X1 Check1_CheckInst_1_U37 ( .A(Red_SignaltoCheck[106]), .B(
        Red_StateRegOutput[46]), .Z(Check1_CheckInst_1_n31) );
  XOR2_X1 Check1_CheckInst_1_U36 ( .A(Red_SignaltoCheck[13]), .B(Red_final[13]), .Z(Check1_CheckInst_1_n32) );
  NOR4_X1 Check1_CheckInst_1_U35 ( .A1(Check1_CheckInst_1_n28), .A2(
        Check1_CheckInst_1_n27), .A3(Check1_CheckInst_1_n26), .A4(
        Check1_CheckInst_1_n25), .ZN(Check1_CheckInst_1_n44) );
  XOR2_X1 Check1_CheckInst_1_U34 ( .A(Red_sel_Key[1]), .B(
        Red_SignaltoCheck[118]), .Z(Check1_CheckInst_1_n25) );
  XOR2_X1 Check1_CheckInst_1_U33 ( .A(Red_RoundConstant[4]), .B(
        Red_SignaltoCheck[112]), .Z(Check1_CheckInst_1_n26) );
  XOR2_X1 Check1_CheckInst_1_U32 ( .A(Red_final[1]), .B(Red_SignaltoCheck[1]), 
        .Z(Check1_CheckInst_1_n27) );
  XOR2_X1 Check1_CheckInst_1_U31 ( .A(Red_StateRegOutput[43]), .B(
        Red_SignaltoCheck[103]), .Z(Check1_CheckInst_1_n28) );
  NAND4_X1 Check1_CheckInst_1_U30 ( .A1(Check1_CheckInst_1_n24), .A2(
        Check1_CheckInst_1_n23), .A3(Check1_CheckInst_1_n22), .A4(
        Check1_CheckInst_1_n21), .ZN(Check1_CheckInst_1_n46) );
  XNOR2_X1 Check1_CheckInst_1_U29 ( .A(Red_final[10]), .B(
        Red_SignaltoCheck[10]), .ZN(Check1_CheckInst_1_n21) );
  XNOR2_X1 Check1_CheckInst_1_U28 ( .A(Red_StateRegOutput[16]), .B(
        Red_SignaltoCheck[76]), .ZN(Check1_CheckInst_1_n22) );
  XNOR2_X1 Check1_CheckInst_1_U27 ( .A(Red_RoundConstant[1]), .B(
        Red_SignaltoCheck[109]), .ZN(Check1_CheckInst_1_n23) );
  NOR4_X1 Check1_CheckInst_1_U26 ( .A1(Check1_CheckInst_1_n20), .A2(
        Check1_CheckInst_1_n19), .A3(Check1_CheckInst_1_n18), .A4(
        Check1_CheckInst_1_n17), .ZN(Check1_CheckInst_1_n24) );
  XOR2_X1 Check1_CheckInst_1_U25 ( .A(Red_final[16]), .B(Red_SignaltoCheck[16]), .Z(Check1_CheckInst_1_n17) );
  XOR2_X1 Check1_CheckInst_1_U24 ( .A(Red_StateRegOutput[19]), .B(
        Red_SignaltoCheck[79]), .Z(Check1_CheckInst_1_n18) );
  XOR2_X1 Check1_CheckInst_1_U23 ( .A(Red_StateRegOutput[13]), .B(
        Red_SignaltoCheck[73]), .Z(Check1_CheckInst_1_n19) );
  XOR2_X1 Check1_CheckInst_1_U22 ( .A(Red_StateRegOutput[28]), .B(
        Red_SignaltoCheck[88]), .Z(Check1_CheckInst_1_n20) );
  XOR2_X1 Check1_CheckInst_1_U21 ( .A(Red_StateRegOutput[4]), .B(
        Red_SignaltoCheck[64]), .Z(Check1_CheckInst_1_n47) );
  XOR2_X1 Check1_CheckInst_1_U20 ( .A(Red_FSMUpdate[1]), .B(
        Red_SignaltoCheck[49]), .Z(Check1_CheckInst_1_n48) );
  NOR3_X1 Check1_CheckInst_1_U19 ( .A1(Check1_CheckInst_1_n16), .A2(
        Check1_CheckInst_1_n15), .A3(Check1_CheckInst_1_n14), .ZN(
        Check1_CheckInst_1_n52) );
  NAND4_X1 Check1_CheckInst_1_U18 ( .A1(Check1_CheckInst_1_n13), .A2(
        Check1_CheckInst_1_n12), .A3(Check1_CheckInst_1_n11), .A4(
        Check1_CheckInst_1_n10), .ZN(Check1_CheckInst_1_n14) );
  XNOR2_X1 Check1_CheckInst_1_U17 ( .A(Red_selectsNext[4]), .B(
        Red_SignaltoCheck[58]), .ZN(Check1_CheckInst_1_n10) );
  XNOR2_X1 Check1_CheckInst_1_U16 ( .A(Red_StateRegOutput[25]), .B(
        Red_SignaltoCheck[85]), .ZN(Check1_CheckInst_1_n11) );
  XNOR2_X1 Check1_CheckInst_1_U15 ( .A(Red_StateRegOutput[10]), .B(
        Red_SignaltoCheck[70]), .ZN(Check1_CheckInst_1_n12) );
  XNOR2_X1 Check1_CheckInst_1_U14 ( .A(Red_StateRegOutput[22]), .B(
        Red_SignaltoCheck[82]), .ZN(Check1_CheckInst_1_n13) );
  XOR2_X1 Check1_CheckInst_1_U13 ( .A(Red_final[4]), .B(Red_SignaltoCheck[4]), 
        .Z(Check1_CheckInst_1_n15) );
  XOR2_X1 Check1_CheckInst_1_U12 ( .A(Red_SignaltoCheck[7]), .B(Red_final[7]), 
        .Z(Check1_CheckInst_1_n16) );
  XNOR2_X1 Check1_CheckInst_1_U11 ( .A(Red_StateRegOutput[1]), .B(
        Red_SignaltoCheck[61]), .ZN(Check1_CheckInst_1_n7) );
  XNOR2_X1 Check1_CheckInst_1_U10 ( .A(Red_SignaltoCheck[67]), .B(
        Red_StateRegOutput[7]), .ZN(Check1_CheckInst_1_n8) );
  NOR4_X1 Check1_CheckInst_1_U9 ( .A1(Check1_CheckInst_1_n6), .A2(
        Check1_CheckInst_1_n5), .A3(Check1_CheckInst_1_n4), .A4(
        Check1_CheckInst_1_n3), .ZN(Check1_CheckInst_1_n9) );
  XOR2_X1 Check1_CheckInst_1_U8 ( .A(Red_StateRegOutput[34]), .B(
        Red_SignaltoCheck[94]), .Z(Check1_CheckInst_1_n3) );
  XOR2_X1 Check1_CheckInst_1_U7 ( .A(Red_StateRegOutput[40]), .B(
        Red_SignaltoCheck[100]), .Z(Check1_CheckInst_1_n4) );
  XOR2_X1 Check1_CheckInst_1_U6 ( .A(Red_selectsNext[1]), .B(
        Red_SignaltoCheck[55]), .Z(Check1_CheckInst_1_n5) );
  XOR2_X1 Check1_CheckInst_1_U5 ( .A(Red_StateRegOutput[31]), .B(
        Red_SignaltoCheck[91]), .Z(Check1_CheckInst_1_n6) );
  XOR2_X1 Check1_CheckInst_1_U4 ( .A(Red_final[46]), .B(Red_SignaltoCheck[46]), 
        .Z(Check1_CheckInst_1_n54) );
  NOR3_X1 Check1_CheckInst_1_U3 ( .A1(Check1_CheckInst_1_n54), .A2(
        Check1_CheckInst_1_n53), .A3(Check1_CheckInst_1_n2), .ZN(Error[1]) );
  NAND4_X1 Check1_CheckInst_1_U2 ( .A1(Check1_CheckInst_1_n9), .A2(
        Check1_CheckInst_1_n7), .A3(Check1_CheckInst_1_n8), .A4(
        Check1_CheckInst_1_n1), .ZN(Check1_CheckInst_1_n2) );
  XNOR2_X1 Check1_CheckInst_1_U1 ( .A(Red_FSMUpdate[4]), .B(
        Red_SignaltoCheck[52]), .ZN(Check1_CheckInst_1_n1) );
  NAND4_X1 Check1_CheckInst_2_U55 ( .A1(Check1_CheckInst_2_n50), .A2(
        Check1_CheckInst_2_n49), .A3(Check1_CheckInst_2_n48), .A4(
        Check1_CheckInst_2_n47), .ZN(Check1_CheckInst_2_n51) );
  XNOR2_X1 Check1_CheckInst_2_U54 ( .A(Red_StateRegOutput[38]), .B(
        Red_SignaltoCheck[98]), .ZN(Check1_CheckInst_2_n47) );
  XNOR2_X1 Check1_CheckInst_2_U53 ( .A(1'b0), .B(Red_SignaltoCheck[122]), .ZN(
        Check1_CheckInst_2_n48) );
  NOR4_X1 Check1_CheckInst_2_U52 ( .A1(Check1_CheckInst_2_n46), .A2(
        Check1_CheckInst_2_n45), .A3(Check1_CheckInst_2_n44), .A4(
        Check1_CheckInst_2_n43), .ZN(Check1_CheckInst_2_n49) );
  NAND4_X1 Check1_CheckInst_2_U51 ( .A1(Check1_CheckInst_2_n42), .A2(
        Check1_CheckInst_2_n41), .A3(Check1_CheckInst_2_n40), .A4(
        Check1_CheckInst_2_n39), .ZN(Check1_CheckInst_2_n43) );
  NOR4_X1 Check1_CheckInst_2_U50 ( .A1(Check1_CheckInst_2_n38), .A2(
        Check1_CheckInst_2_n37), .A3(Check1_CheckInst_2_n36), .A4(
        Check1_CheckInst_2_n35), .ZN(Check1_CheckInst_2_n39) );
  XOR2_X1 Check1_CheckInst_2_U49 ( .A(Red_final[44]), .B(Red_SignaltoCheck[44]), .Z(Check1_CheckInst_2_n35) );
  XOR2_X1 Check1_CheckInst_2_U48 ( .A(Red_final[35]), .B(Red_SignaltoCheck[35]), .Z(Check1_CheckInst_2_n36) );
  XOR2_X1 Check1_CheckInst_2_U47 ( .A(Red_final[41]), .B(Red_SignaltoCheck[41]), .Z(Check1_CheckInst_2_n37) );
  XOR2_X1 Check1_CheckInst_2_U46 ( .A(Red_final[38]), .B(Red_SignaltoCheck[38]), .Z(Check1_CheckInst_2_n38) );
  NOR4_X1 Check1_CheckInst_2_U45 ( .A1(Check1_CheckInst_2_n34), .A2(
        Check1_CheckInst_2_n33), .A3(Check1_CheckInst_2_n32), .A4(
        Check1_CheckInst_2_n31), .ZN(Check1_CheckInst_2_n40) );
  XOR2_X1 Check1_CheckInst_2_U44 ( .A(Red_final[32]), .B(Red_SignaltoCheck[32]), .Z(Check1_CheckInst_2_n31) );
  XOR2_X1 Check1_CheckInst_2_U43 ( .A(Red_final[29]), .B(Red_SignaltoCheck[29]), .Z(Check1_CheckInst_2_n32) );
  XOR2_X1 Check1_CheckInst_2_U42 ( .A(Red_final[20]), .B(Red_SignaltoCheck[20]), .Z(Check1_CheckInst_2_n33) );
  XOR2_X1 Check1_CheckInst_2_U41 ( .A(Red_final[26]), .B(Red_SignaltoCheck[26]), .Z(Check1_CheckInst_2_n34) );
  NOR4_X1 Check1_CheckInst_2_U40 ( .A1(Check1_CheckInst_2_n30), .A2(
        Check1_CheckInst_2_n29), .A3(Check1_CheckInst_2_n28), .A4(
        Check1_CheckInst_2_n27), .ZN(Check1_CheckInst_2_n41) );
  XOR2_X1 Check1_CheckInst_2_U39 ( .A(Red_final[23]), .B(Red_SignaltoCheck[23]), .Z(Check1_CheckInst_2_n27) );
  XOR2_X1 Check1_CheckInst_2_U38 ( .A(Red_sel_Tweak[2]), .B(
        Red_SignaltoCheck[116]), .Z(Check1_CheckInst_2_n28) );
  XOR2_X1 Check1_CheckInst_2_U37 ( .A(Red_SignaltoCheck[107]), .B(
        Red_StateRegOutput[47]), .Z(Check1_CheckInst_2_n29) );
  XOR2_X1 Check1_CheckInst_2_U36 ( .A(Red_SignaltoCheck[14]), .B(Red_final[14]), .Z(Check1_CheckInst_2_n30) );
  NOR4_X1 Check1_CheckInst_2_U35 ( .A1(Check1_CheckInst_2_n26), .A2(
        Check1_CheckInst_2_n25), .A3(Check1_CheckInst_2_n24), .A4(
        Check1_CheckInst_2_n23), .ZN(Check1_CheckInst_2_n42) );
  XOR2_X1 Check1_CheckInst_2_U34 ( .A(Red_sel_Key[2]), .B(
        Red_SignaltoCheck[119]), .Z(Check1_CheckInst_2_n23) );
  XOR2_X1 Check1_CheckInst_2_U33 ( .A(Red_RoundConstant[5]), .B(
        Red_SignaltoCheck[113]), .Z(Check1_CheckInst_2_n24) );
  XOR2_X1 Check1_CheckInst_2_U32 ( .A(Red_final[2]), .B(Red_SignaltoCheck[2]), 
        .Z(Check1_CheckInst_2_n25) );
  XOR2_X1 Check1_CheckInst_2_U31 ( .A(Red_StateRegOutput[44]), .B(
        Red_SignaltoCheck[104]), .Z(Check1_CheckInst_2_n26) );
  NAND4_X1 Check1_CheckInst_2_U30 ( .A1(Check1_CheckInst_2_n22), .A2(
        Check1_CheckInst_2_n21), .A3(Check1_CheckInst_2_n20), .A4(
        Check1_CheckInst_2_n19), .ZN(Check1_CheckInst_2_n44) );
  XNOR2_X1 Check1_CheckInst_2_U29 ( .A(Red_final[11]), .B(
        Red_SignaltoCheck[11]), .ZN(Check1_CheckInst_2_n19) );
  XNOR2_X1 Check1_CheckInst_2_U28 ( .A(Red_StateRegOutput[17]), .B(
        Red_SignaltoCheck[77]), .ZN(Check1_CheckInst_2_n20) );
  XNOR2_X1 Check1_CheckInst_2_U27 ( .A(Red_RoundConstant[2]), .B(
        Red_SignaltoCheck[110]), .ZN(Check1_CheckInst_2_n21) );
  NOR4_X1 Check1_CheckInst_2_U26 ( .A1(Check1_CheckInst_2_n18), .A2(
        Check1_CheckInst_2_n17), .A3(Check1_CheckInst_2_n16), .A4(
        Check1_CheckInst_2_n15), .ZN(Check1_CheckInst_2_n22) );
  XOR2_X1 Check1_CheckInst_2_U25 ( .A(Red_final[17]), .B(Red_SignaltoCheck[17]), .Z(Check1_CheckInst_2_n15) );
  XOR2_X1 Check1_CheckInst_2_U24 ( .A(Red_StateRegOutput[20]), .B(
        Red_SignaltoCheck[80]), .Z(Check1_CheckInst_2_n16) );
  XOR2_X1 Check1_CheckInst_2_U23 ( .A(Red_StateRegOutput[14]), .B(
        Red_SignaltoCheck[74]), .Z(Check1_CheckInst_2_n17) );
  XOR2_X1 Check1_CheckInst_2_U22 ( .A(Red_StateRegOutput[29]), .B(
        Red_SignaltoCheck[89]), .Z(Check1_CheckInst_2_n18) );
  XOR2_X1 Check1_CheckInst_2_U21 ( .A(Red_StateRegOutput[5]), .B(
        Red_SignaltoCheck[65]), .Z(Check1_CheckInst_2_n45) );
  XOR2_X1 Check1_CheckInst_2_U20 ( .A(Red_FSMUpdate[2]), .B(
        Red_SignaltoCheck[50]), .Z(Check1_CheckInst_2_n46) );
  NOR3_X1 Check1_CheckInst_2_U19 ( .A1(Check1_CheckInst_2_n14), .A2(
        Check1_CheckInst_2_n13), .A3(Check1_CheckInst_2_n12), .ZN(
        Check1_CheckInst_2_n50) );
  NAND4_X1 Check1_CheckInst_2_U18 ( .A1(Check1_CheckInst_2_n11), .A2(
        Check1_CheckInst_2_n10), .A3(Check1_CheckInst_2_n9), .A4(
        Check1_CheckInst_2_n8), .ZN(Check1_CheckInst_2_n12) );
  XNOR2_X1 Check1_CheckInst_2_U17 ( .A(1'b0), .B(Red_SignaltoCheck[59]), .ZN(
        Check1_CheckInst_2_n8) );
  XNOR2_X1 Check1_CheckInst_2_U16 ( .A(Red_StateRegOutput[26]), .B(
        Red_SignaltoCheck[86]), .ZN(Check1_CheckInst_2_n9) );
  XNOR2_X1 Check1_CheckInst_2_U15 ( .A(Red_StateRegOutput[11]), .B(
        Red_SignaltoCheck[71]), .ZN(Check1_CheckInst_2_n10) );
  XNOR2_X1 Check1_CheckInst_2_U14 ( .A(Red_StateRegOutput[23]), .B(
        Red_SignaltoCheck[83]), .ZN(Check1_CheckInst_2_n11) );
  XOR2_X1 Check1_CheckInst_2_U13 ( .A(Red_final[5]), .B(Red_SignaltoCheck[5]), 
        .Z(Check1_CheckInst_2_n13) );
  XOR2_X1 Check1_CheckInst_2_U12 ( .A(Red_SignaltoCheck[8]), .B(Red_final[8]), 
        .Z(Check1_CheckInst_2_n14) );
  NAND3_X1 Check1_CheckInst_2_U11 ( .A1(Check1_CheckInst_2_n7), .A2(
        Check1_CheckInst_2_n6), .A3(Check1_CheckInst_2_n5), .ZN(
        Check1_CheckInst_2_n52) );
  XNOR2_X1 Check1_CheckInst_2_U10 ( .A(Red_StateRegOutput[2]), .B(
        Red_SignaltoCheck[62]), .ZN(Check1_CheckInst_2_n5) );
  XNOR2_X1 Check1_CheckInst_2_U9 ( .A(Red_SignaltoCheck[68]), .B(
        Red_StateRegOutput[8]), .ZN(Check1_CheckInst_2_n6) );
  NOR4_X1 Check1_CheckInst_2_U8 ( .A1(Check1_CheckInst_2_n4), .A2(
        Check1_CheckInst_2_n3), .A3(Check1_CheckInst_2_n2), .A4(
        Check1_CheckInst_2_n1), .ZN(Check1_CheckInst_2_n7) );
  XOR2_X1 Check1_CheckInst_2_U7 ( .A(Red_StateRegOutput[35]), .B(
        Red_SignaltoCheck[95]), .Z(Check1_CheckInst_2_n1) );
  XOR2_X1 Check1_CheckInst_2_U6 ( .A(Red_StateRegOutput[41]), .B(
        Red_SignaltoCheck[101]), .Z(Check1_CheckInst_2_n2) );
  XOR2_X1 Check1_CheckInst_2_U5 ( .A(1'b0), .B(Red_SignaltoCheck[56]), .Z(
        Check1_CheckInst_2_n3) );
  XOR2_X1 Check1_CheckInst_2_U4 ( .A(Red_StateRegOutput[32]), .B(
        Red_SignaltoCheck[92]), .Z(Check1_CheckInst_2_n4) );
  XOR2_X1 Check1_CheckInst_2_U3 ( .A(Red_FSMUpdate[5]), .B(
        Red_SignaltoCheck[53]), .Z(Check1_CheckInst_2_n53) );
  XOR2_X1 Check1_CheckInst_2_U2 ( .A(Red_final[47]), .B(Red_SignaltoCheck[47]), 
        .Z(Check1_CheckInst_2_n54) );
  NOR4_X2 Check1_CheckInst_2_U1 ( .A1(Check1_CheckInst_2_n54), .A2(
        Check1_CheckInst_2_n53), .A3(Check1_CheckInst_2_n52), .A4(
        Check1_CheckInst_2_n51), .ZN(Error[2]) );
  NOR2_X1 ANDInst_0_U3 ( .A1(ANDInst_0_n2), .A2(ANDInst_0_n1), .ZN(
        ErrorFreeUpdate[0]) );
  NAND4_X1 ANDInst_0_U2 ( .A1(ErrorFree[2]), .A2(ErrorFree[3]), .A3(
        ErrorFree[0]), .A4(ErrorFree[1]), .ZN(ANDInst_0_n1) );
  NAND4_X1 ANDInst_0_U1 ( .A1(Error[1]), .A2(Error[2]), .A3(ErrorFree[4]), 
        .A4(Error[0]), .ZN(ANDInst_0_n2) );
  NOR2_X1 ANDInst_1_U3 ( .A1(ANDInst_1_n2), .A2(ANDInst_1_n1), .ZN(
        ErrorFreeUpdate[1]) );
  NAND4_X1 ANDInst_1_U2 ( .A1(ErrorFree[2]), .A2(ErrorFree[3]), .A3(
        ErrorFree[0]), .A4(ErrorFree[1]), .ZN(ANDInst_1_n1) );
  NAND4_X1 ANDInst_1_U1 ( .A1(Error[1]), .A2(Error[2]), .A3(ErrorFree[4]), 
        .A4(Error[0]), .ZN(ANDInst_1_n2) );
  NOR2_X1 ANDInst_2_U3 ( .A1(ANDInst_2_n2), .A2(ANDInst_2_n1), .ZN(
        ErrorFreeUpdate[2]) );
  NAND4_X1 ANDInst_2_U2 ( .A1(ErrorFree[2]), .A2(ErrorFree[3]), .A3(
        ErrorFree[0]), .A4(ErrorFree[1]), .ZN(ANDInst_2_n1) );
  NAND4_X1 ANDInst_2_U1 ( .A1(Error[1]), .A2(Error[2]), .A3(ErrorFree[4]), 
        .A4(Error[0]), .ZN(ANDInst_2_n2) );
  NAND4_X1 ANDInst_3_U3 ( .A1(ErrorFree[2]), .A2(ErrorFree[3]), .A3(
        ErrorFree[0]), .A4(ErrorFree[1]), .ZN(ANDInst_3_n1) );
  NAND4_X1 ANDInst_3_U2 ( .A1(Error[1]), .A2(Error[2]), .A3(ErrorFree[4]), 
        .A4(Error[0]), .ZN(ANDInst_3_n2) );
  NOR2_X1 ANDInst_3_U1 ( .A1(ANDInst_3_n2), .A2(ANDInst_3_n1), .ZN(
        ErrorFreeUpdate[3]) );
  NAND4_X1 ANDInst_4_U3 ( .A1(ErrorFree[2]), .A2(ErrorFree[3]), .A3(
        ErrorFree[0]), .A4(ErrorFree[1]), .ZN(ANDInst_4_n1) );
  NAND4_X1 ANDInst_4_U2 ( .A1(Error[1]), .A2(Error[2]), .A3(ErrorFree[4]), 
        .A4(Error[0]), .ZN(ANDInst_4_n2) );
  NOR2_X1 ANDInst_4_U1 ( .A1(ANDInst_4_n2), .A2(ANDInst_4_n1), .ZN(
        ErrorFreeUpdate[4]) );
  BUF_X1 OutputMUX_U15 ( .A(ErrorFreeUpdate[0]), .Z(OutputMUX_n2) );
  BUF_X1 OutputMUX_U14 ( .A(ErrorFreeUpdate[0]), .Z(OutputMUX_n1) );
  BUF_X1 OutputMUX_U13 ( .A(ErrorFreeUpdate[1]), .Z(OutputMUX_n5) );
  BUF_X1 OutputMUX_U12 ( .A(OutputMUX_n1), .Z(OutputMUX_n3) );
  BUF_X1 OutputMUX_U11 ( .A(ErrorFreeUpdate[2]), .Z(OutputMUX_n8) );
  BUF_X1 OutputMUX_U10 ( .A(ErrorFreeUpdate[3]), .Z(OutputMUX_n11) );
  BUF_X1 OutputMUX_U9 ( .A(ErrorFreeUpdate[4]), .Z(OutputMUX_n14) );
  BUF_X1 OutputMUX_U8 ( .A(ErrorFreeUpdate[1]), .Z(OutputMUX_n4) );
  BUF_X1 OutputMUX_U7 ( .A(ErrorFreeUpdate[2]), .Z(OutputMUX_n7) );
  BUF_X1 OutputMUX_U6 ( .A(OutputMUX_n4), .Z(OutputMUX_n6) );
  BUF_X1 OutputMUX_U5 ( .A(OutputMUX_n7), .Z(OutputMUX_n9) );
  BUF_X1 OutputMUX_U4 ( .A(OutputMUX_n10), .Z(OutputMUX_n12) );
  BUF_X1 OutputMUX_U3 ( .A(ErrorFreeUpdate[3]), .Z(OutputMUX_n10) );
  BUF_X1 OutputMUX_U2 ( .A(ErrorFreeUpdate[4]), .Z(OutputMUX_n13) );
  BUF_X1 OutputMUX_U1 ( .A(OutputMUX_n13), .Z(OutputMUX_n15) );
  MUX2_X1 OutputMUX_MUX2to1Inst_0_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[60]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_0_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_0_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_0_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_0_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_0_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_0_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_0_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_0_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_0_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_0_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_0_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_0_sig[4]), .S(OutputMUX_n15), .Z(OutputRegIn[0])
         );
  MUX2_X1 OutputMUX_MUX2to1Inst_1_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[61]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_1_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_1_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_1_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_1_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_1_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_1_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_1_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_1_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_1_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_1_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_1_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_1_sig[4]), .S(OutputMUX_n14), .Z(OutputRegIn[1])
         );
  MUX2_X1 OutputMUX_MUX2to1Inst_2_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[62]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_2_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_2_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_2_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_2_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_2_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_2_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_2_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_2_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_2_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_2_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_2_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_2_sig[4]), .S(OutputMUX_n14), .Z(OutputRegIn[2])
         );
  MUX2_X1 OutputMUX_MUX2to1Inst_3_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[63]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_3_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_3_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_3_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_3_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_3_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_3_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_3_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_3_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_3_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_3_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_3_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_3_sig[4]), .S(OutputMUX_n14), .Z(OutputRegIn[3])
         );
  MUX2_X1 OutputMUX_MUX2to1Inst_4_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[48]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_4_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_4_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_4_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_4_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_4_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_4_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_4_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_4_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_4_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_4_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_4_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_4_sig[4]), .S(OutputMUX_n14), .Z(OutputRegIn[4])
         );
  MUX2_X1 OutputMUX_MUX2to1Inst_5_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[49]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_5_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_5_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_5_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_5_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_5_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_5_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_5_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_5_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_5_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_5_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_5_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_5_sig[4]), .S(OutputMUX_n14), .Z(OutputRegIn[5])
         );
  MUX2_X1 OutputMUX_MUX2to1Inst_6_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[50]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_6_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_6_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_6_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_6_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_6_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_6_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_6_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_6_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_6_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_6_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_6_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_6_sig[4]), .S(OutputMUX_n14), .Z(OutputRegIn[6])
         );
  MUX2_X1 OutputMUX_MUX2to1Inst_7_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[51]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_7_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_7_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_7_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_7_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_7_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_7_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_7_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_7_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_7_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_7_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_7_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_7_sig[4]), .S(OutputMUX_n14), .Z(OutputRegIn[7])
         );
  MUX2_X1 OutputMUX_MUX2to1Inst_8_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[52]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_8_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_8_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_8_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_8_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_8_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_8_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_8_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_8_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_8_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_8_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_8_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_8_sig[4]), .S(OutputMUX_n14), .Z(OutputRegIn[8])
         );
  MUX2_X1 OutputMUX_MUX2to1Inst_9_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[53]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_9_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_9_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_9_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_9_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_9_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_9_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_9_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_9_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_9_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_9_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_9_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_9_sig[4]), .S(OutputMUX_n14), .Z(OutputRegIn[9])
         );
  MUX2_X1 OutputMUX_MUX2to1Inst_10_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[54]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_10_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_10_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_10_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_10_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_10_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_10_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_10_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_10_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_10_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_10_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_10_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_10_sig[4]), .S(OutputMUX_n14), .Z(
        OutputRegIn[10]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_11_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[55]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_11_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_11_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_11_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_11_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_11_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_11_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_11_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_11_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_11_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_11_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_11_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_11_sig[4]), .S(OutputMUX_n14), .Z(
        OutputRegIn[11]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_12_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[56]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_12_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_12_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_12_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_12_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_12_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_12_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_12_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_12_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_12_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_12_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_12_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_12_sig[4]), .S(OutputMUX_n14), .Z(
        OutputRegIn[12]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_13_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[57]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_13_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_13_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_13_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_13_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_13_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_13_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_13_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_13_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_13_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_13_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_13_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_13_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[13]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_14_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[58]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_14_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_14_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_14_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_14_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_14_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_14_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_14_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_14_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_14_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_14_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_14_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_14_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[14]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_15_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[59]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_15_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_15_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_15_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_15_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_15_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_15_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_15_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_15_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_15_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_15_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_15_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_15_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[15]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_16_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[32]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_16_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_16_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_16_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_16_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_16_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_16_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_16_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_16_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_16_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_16_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_16_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_16_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[16]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_17_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[33]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_17_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_17_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_17_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_17_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_17_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_17_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_17_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_17_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_17_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_17_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_17_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_17_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[17]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_18_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[34]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_18_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_18_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_18_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_18_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_18_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_18_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_18_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_18_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_18_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_18_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_18_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_18_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[18]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_19_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[35]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_19_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_19_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_19_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_19_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_19_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_19_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_19_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_19_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_19_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_19_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_19_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_19_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[19]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_20_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[44]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_20_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_20_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_20_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_20_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_20_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_20_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_20_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_20_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_20_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_20_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_20_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_20_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[20]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_21_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[45]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_21_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_21_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_21_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_21_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_21_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_21_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_21_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_21_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_21_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_21_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_21_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_21_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[21]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_22_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[46]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_22_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_22_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_22_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_22_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_22_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_22_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_22_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_22_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_22_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_22_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_22_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_22_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[22]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_23_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[47]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_23_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_23_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_23_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_23_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_23_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_23_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_23_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_23_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_23_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_23_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_23_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_23_sig[4]), .S(OutputMUX_n14), .Z(
        OutputRegIn[23]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_24_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[40]), .S(OutputMUX_n1), .Z(
        OutputMUX_MUX2to1Inst_24_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_24_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_24_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_24_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_24_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_24_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_24_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_24_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_24_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_24_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_24_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_24_sig[4]), .S(OutputMUX_n14), .Z(
        OutputRegIn[24]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_25_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[41]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_25_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_25_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_25_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_25_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_25_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_25_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_25_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_25_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_25_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_25_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_25_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_25_sig[4]), .S(OutputMUX_n14), .Z(
        OutputRegIn[25]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_26_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[42]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_26_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_26_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_26_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_26_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_26_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_26_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_26_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_26_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_26_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_26_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_26_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_26_sig[4]), .S(OutputMUX_n14), .Z(
        OutputRegIn[26]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_27_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[43]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_27_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_27_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_27_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_27_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_27_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_27_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_27_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_27_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_27_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_27_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_27_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_27_sig[4]), .S(OutputMUX_n14), .Z(
        OutputRegIn[27]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_28_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[36]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_28_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_28_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_28_sig[1]), .S(OutputMUX_n5), .Z(
        OutputMUX_MUX2to1Inst_28_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_28_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_28_sig[2]), .S(OutputMUX_n8), .Z(
        OutputMUX_MUX2to1Inst_28_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_28_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_28_sig[3]), .S(OutputMUX_n11), .Z(
        OutputMUX_MUX2to1Inst_28_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_28_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_28_sig[4]), .S(OutputMUX_n14), .Z(
        OutputRegIn[28]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_29_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[37]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_29_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_29_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_29_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_29_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_29_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_29_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_29_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_29_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_29_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_29_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_29_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_29_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[29]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_30_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[38]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_30_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_30_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_30_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_30_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_30_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_30_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_30_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_30_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_30_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_30_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_30_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_30_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[30]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_31_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[39]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_31_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_31_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_31_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_31_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_31_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_31_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_31_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_31_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_31_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_31_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_31_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_31_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[31]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_32_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[16]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_32_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_32_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_32_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_32_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_32_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_32_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_32_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_32_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_32_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_32_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_32_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_32_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[32]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_33_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[17]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_33_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_33_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_33_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_33_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_33_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_33_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_33_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_33_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_33_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_33_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_33_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_33_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[33]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_34_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[18]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_34_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_34_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_34_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_34_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_34_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_34_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_34_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_34_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_34_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_34_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_34_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_34_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[34]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_35_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[19]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_35_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_35_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_35_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_35_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_35_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_35_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_35_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_35_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_35_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_35_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_35_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_35_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[35]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_36_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[28]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_36_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_36_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_36_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_36_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_36_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_36_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_36_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_36_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_36_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_36_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_36_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_36_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[36]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_37_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[29]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_37_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_37_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_37_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_37_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_37_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_37_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_37_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_37_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_37_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_37_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_37_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_37_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[37]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_38_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[30]), .S(ErrorFreeUpdate[0]), .Z(
        OutputMUX_MUX2to1Inst_38_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_38_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_38_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_38_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_38_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_38_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_38_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_38_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_38_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_38_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_38_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_38_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[38]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_39_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[31]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_39_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_39_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_39_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_39_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_39_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_39_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_39_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_39_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_39_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_39_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_39_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_39_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[39]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_40_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[24]), .S(ErrorFreeUpdate[0]), .Z(
        OutputMUX_MUX2to1Inst_40_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_40_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_40_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_40_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_40_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_40_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_40_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_40_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_40_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_40_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_40_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_40_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[40]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_41_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[25]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_41_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_41_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_41_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_41_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_41_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_41_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_41_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_41_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_41_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_41_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_41_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_41_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[41]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_42_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[26]), .S(ErrorFreeUpdate[0]), .Z(
        OutputMUX_MUX2to1Inst_42_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_42_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_42_sig[1]), .S(ErrorFreeUpdate[1]), .Z(
        OutputMUX_MUX2to1Inst_42_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_42_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_42_sig[2]), .S(ErrorFreeUpdate[2]), .Z(
        OutputMUX_MUX2to1Inst_42_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_42_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_42_sig[3]), .S(ErrorFreeUpdate[3]), .Z(
        OutputMUX_MUX2to1Inst_42_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_42_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_42_sig[4]), .S(ErrorFreeUpdate[4]), .Z(
        OutputRegIn[42]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_43_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[27]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_43_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_43_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_43_sig[1]), .S(ErrorFreeUpdate[1]), .Z(
        OutputMUX_MUX2to1Inst_43_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_43_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_43_sig[2]), .S(ErrorFreeUpdate[2]), .Z(
        OutputMUX_MUX2to1Inst_43_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_43_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_43_sig[3]), .S(ErrorFreeUpdate[3]), .Z(
        OutputMUX_MUX2to1Inst_43_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_43_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_43_sig[4]), .S(ErrorFreeUpdate[4]), .Z(
        OutputRegIn[43]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_44_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[20]), .S(ErrorFreeUpdate[0]), .Z(
        OutputMUX_MUX2to1Inst_44_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_44_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_44_sig[1]), .S(ErrorFreeUpdate[1]), .Z(
        OutputMUX_MUX2to1Inst_44_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_44_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_44_sig[2]), .S(ErrorFreeUpdate[2]), .Z(
        OutputMUX_MUX2to1Inst_44_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_44_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_44_sig[3]), .S(ErrorFreeUpdate[3]), .Z(
        OutputMUX_MUX2to1Inst_44_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_44_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_44_sig[4]), .S(ErrorFreeUpdate[4]), .Z(
        OutputRegIn[44]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_45_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[21]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_45_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_45_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_45_sig[1]), .S(ErrorFreeUpdate[1]), .Z(
        OutputMUX_MUX2to1Inst_45_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_45_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_45_sig[2]), .S(ErrorFreeUpdate[2]), .Z(
        OutputMUX_MUX2to1Inst_45_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_45_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_45_sig[3]), .S(ErrorFreeUpdate[3]), .Z(
        OutputMUX_MUX2to1Inst_45_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_45_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_45_sig[4]), .S(ErrorFreeUpdate[4]), .Z(
        OutputRegIn[45]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_46_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[22]), .S(ErrorFreeUpdate[0]), .Z(
        OutputMUX_MUX2to1Inst_46_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_46_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_46_sig[1]), .S(ErrorFreeUpdate[1]), .Z(
        OutputMUX_MUX2to1Inst_46_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_46_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_46_sig[2]), .S(ErrorFreeUpdate[2]), .Z(
        OutputMUX_MUX2to1Inst_46_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_46_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_46_sig[3]), .S(ErrorFreeUpdate[3]), .Z(
        OutputMUX_MUX2to1Inst_46_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_46_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_46_sig[4]), .S(ErrorFreeUpdate[4]), .Z(
        OutputRegIn[46]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_47_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[23]), .S(ErrorFreeUpdate[0]), .Z(
        OutputMUX_MUX2to1Inst_47_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_47_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_47_sig[1]), .S(ErrorFreeUpdate[1]), .Z(
        OutputMUX_MUX2to1Inst_47_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_47_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_47_sig[2]), .S(ErrorFreeUpdate[2]), .Z(
        OutputMUX_MUX2to1Inst_47_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_47_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_47_sig[3]), .S(ErrorFreeUpdate[3]), .Z(
        OutputMUX_MUX2to1Inst_47_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_47_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_47_sig[4]), .S(ErrorFreeUpdate[4]), .Z(
        OutputRegIn[47]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_48_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[4]), .S(ErrorFreeUpdate[0]), .Z(
        OutputMUX_MUX2to1Inst_48_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_48_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_48_sig[1]), .S(ErrorFreeUpdate[1]), .Z(
        OutputMUX_MUX2to1Inst_48_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_48_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_48_sig[2]), .S(ErrorFreeUpdate[2]), .Z(
        OutputMUX_MUX2to1Inst_48_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_48_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_48_sig[3]), .S(ErrorFreeUpdate[3]), .Z(
        OutputMUX_MUX2to1Inst_48_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_48_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_48_sig[4]), .S(ErrorFreeUpdate[4]), .Z(
        OutputRegIn[48]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_49_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[5]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_49_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_49_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_49_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_49_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_49_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_49_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_49_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_49_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_49_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_49_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_49_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_49_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[49]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_50_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[6]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_50_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_50_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_50_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_50_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_50_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_50_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_50_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_50_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_50_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_50_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_50_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_50_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[50]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_51_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[7]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_51_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_51_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_51_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_51_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_51_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_51_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_51_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_51_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_51_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_51_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_51_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_51_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[51]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_52_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[8]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_52_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_52_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_52_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_52_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_52_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_52_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_52_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_52_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_52_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_52_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_52_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_52_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[52]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_53_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[9]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_53_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_53_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_53_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_53_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_53_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_53_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_53_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_53_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_53_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_53_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_53_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_53_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[53]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_54_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[10]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_54_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_54_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_54_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_54_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_54_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_54_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_54_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_54_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_54_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_54_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_54_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_54_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[54]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_55_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[11]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_55_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_55_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_55_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_55_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_55_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_55_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_55_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_55_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_55_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_55_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_55_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_55_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[55]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_56_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[12]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_56_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_56_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_56_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_56_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_56_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_56_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_56_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_56_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_56_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_56_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_56_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_56_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[56]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_57_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[13]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_57_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_57_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_57_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_57_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_57_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_57_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_57_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_57_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_57_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_57_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_57_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_57_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[57]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_58_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[14]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_58_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_58_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_58_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_58_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_58_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_58_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_58_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_58_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_58_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_58_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_58_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_58_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[58]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_59_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[15]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_59_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_59_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_59_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_59_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_59_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_59_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_59_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_59_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_59_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_59_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_59_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_59_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[59]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_60_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[0]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_60_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_60_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_60_sig[1]), .S(OutputMUX_n6), .Z(
        OutputMUX_MUX2to1Inst_60_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_60_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_60_sig[2]), .S(OutputMUX_n9), .Z(
        OutputMUX_MUX2to1Inst_60_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_60_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_60_sig[3]), .S(OutputMUX_n12), .Z(
        OutputMUX_MUX2to1Inst_60_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_60_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_60_sig[4]), .S(OutputMUX_n15), .Z(
        OutputRegIn[60]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_61_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[1]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_61_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_61_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_61_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_61_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_61_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_61_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_61_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_61_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_61_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_61_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_61_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_61_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[61]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_62_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[2]), .S(OutputMUX_n3), .Z(
        OutputMUX_MUX2to1Inst_62_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_62_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_62_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_62_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_62_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_62_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_62_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_62_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_62_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_62_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_62_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_62_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[62]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_63_MUXInst_0_U1 ( .A(1'b0), .B(
        PermutationOutput[3]), .S(OutputMUX_n2), .Z(
        OutputMUX_MUX2to1Inst_63_sig[1]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_63_MUXInst_1_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_63_sig[1]), .S(OutputMUX_n4), .Z(
        OutputMUX_MUX2to1Inst_63_sig[2]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_63_MUXInst_2_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_63_sig[2]), .S(OutputMUX_n7), .Z(
        OutputMUX_MUX2to1Inst_63_sig[3]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_63_MUXInst_3_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_63_sig[3]), .S(OutputMUX_n10), .Z(
        OutputMUX_MUX2to1Inst_63_sig[4]) );
  MUX2_X1 OutputMUX_MUX2to1Inst_63_MUXInst_4_U1 ( .A(1'b0), .B(
        OutputMUX_MUX2to1Inst_63_sig[4]), .S(OutputMUX_n13), .Z(
        OutputRegIn[63]) );
  AOI22_X1 OutputReg_U73 ( .A1(OutputReg_n69), .A2(Output[0]), .B1(
        OutputReg_n2), .B2(OutputRegIn[0]), .ZN(OutputReg_n1) );
  AOI22_X1 OutputReg_U72 ( .A1(OutputReg_n68), .A2(Output[1]), .B1(
        OutputReg_n70), .B2(OutputRegIn[1]), .ZN(OutputReg_n4) );
  AOI22_X1 OutputReg_U71 ( .A1(OutputReg_n68), .A2(Output[2]), .B1(
        OutputReg_n3), .B2(OutputRegIn[2]), .ZN(OutputReg_n5) );
  AOI22_X1 OutputReg_U70 ( .A1(OutputReg_n68), .A2(Output[3]), .B1(
        OutputReg_n2), .B2(OutputRegIn[3]), .ZN(OutputReg_n6) );
  AOI22_X1 OutputReg_U69 ( .A1(OutputReg_n68), .A2(Output[4]), .B1(
        OutputReg_n67), .B2(OutputRegIn[4]), .ZN(OutputReg_n7) );
  AOI22_X1 OutputReg_U68 ( .A1(OutputReg_n68), .A2(Output[5]), .B1(
        OutputReg_n67), .B2(OutputRegIn[5]), .ZN(OutputReg_n8) );
  AOI22_X1 OutputReg_U67 ( .A1(OutputReg_n68), .A2(Output[6]), .B1(
        OutputReg_n67), .B2(OutputRegIn[6]), .ZN(OutputReg_n9) );
  AOI22_X1 OutputReg_U66 ( .A1(OutputReg_n68), .A2(Output[7]), .B1(
        OutputReg_n67), .B2(OutputRegIn[7]), .ZN(OutputReg_n10) );
  AOI22_X1 OutputReg_U65 ( .A1(OutputReg_n68), .A2(Output[8]), .B1(
        OutputReg_n67), .B2(OutputRegIn[8]), .ZN(OutputReg_n11) );
  AOI22_X1 OutputReg_U64 ( .A1(OutputReg_n68), .A2(Output[9]), .B1(
        OutputReg_n67), .B2(OutputRegIn[9]), .ZN(OutputReg_n12) );
  AOI22_X1 OutputReg_U63 ( .A1(OutputReg_n68), .A2(Output[10]), .B1(
        OutputReg_n3), .B2(OutputRegIn[10]), .ZN(OutputReg_n13) );
  AOI22_X1 OutputReg_U62 ( .A1(OutputReg_n69), .A2(Output[11]), .B1(
        OutputReg_n3), .B2(OutputRegIn[11]), .ZN(OutputReg_n14) );
  AOI22_X1 OutputReg_U61 ( .A1(OutputReg_n69), .A2(Output[12]), .B1(
        OutputReg_n2), .B2(OutputRegIn[12]), .ZN(OutputReg_n15) );
  AOI22_X1 OutputReg_U60 ( .A1(OutputReg_n69), .A2(Output[13]), .B1(
        OutputReg_n67), .B2(OutputRegIn[13]), .ZN(OutputReg_n16) );
  AOI22_X1 OutputReg_U59 ( .A1(OutputReg_n69), .A2(Output[14]), .B1(
        OutputReg_n70), .B2(OutputRegIn[14]), .ZN(OutputReg_n17) );
  AOI22_X1 OutputReg_U58 ( .A1(OutputReg_n71), .A2(Output[15]), .B1(
        OutputReg_n70), .B2(OutputRegIn[15]), .ZN(OutputReg_n18) );
  AOI22_X1 OutputReg_U57 ( .A1(OutputReg_n71), .A2(Output[16]), .B1(
        OutputReg_n2), .B2(OutputRegIn[16]), .ZN(OutputReg_n19) );
  AOI22_X1 OutputReg_U56 ( .A1(OutputReg_n69), .A2(Output[17]), .B1(
        OutputReg_n3), .B2(OutputRegIn[17]), .ZN(OutputReg_n20) );
  AOI22_X1 OutputReg_U55 ( .A1(OutputReg_n69), .A2(Output[18]), .B1(
        OutputReg_n2), .B2(OutputRegIn[18]), .ZN(OutputReg_n21) );
  AOI22_X1 OutputReg_U54 ( .A1(OutputReg_n69), .A2(Output[19]), .B1(
        OutputReg_n3), .B2(OutputRegIn[19]), .ZN(OutputReg_n22) );
  AOI22_X1 OutputReg_U53 ( .A1(OutputReg_n69), .A2(Output[20]), .B1(
        OutputReg_n2), .B2(OutputRegIn[20]), .ZN(OutputReg_n23) );
  AOI22_X1 OutputReg_U52 ( .A1(OutputReg_n69), .A2(Output[21]), .B1(
        OutputReg_n3), .B2(OutputRegIn[21]), .ZN(OutputReg_n24) );
  AOI22_X1 OutputReg_U51 ( .A1(OutputReg_n69), .A2(Output[22]), .B1(
        OutputReg_n2), .B2(OutputRegIn[22]), .ZN(OutputReg_n25) );
  AOI22_X1 OutputReg_U50 ( .A1(OutputReg_n69), .A2(Output[23]), .B1(
        OutputReg_n3), .B2(OutputRegIn[23]), .ZN(OutputReg_n26) );
  AOI22_X1 OutputReg_U49 ( .A1(OutputReg_n69), .A2(Output[24]), .B1(
        OutputReg_n2), .B2(OutputRegIn[24]), .ZN(OutputReg_n27) );
  AOI22_X1 OutputReg_U48 ( .A1(OutputReg_n69), .A2(Output[25]), .B1(
        OutputReg_n3), .B2(OutputRegIn[25]), .ZN(OutputReg_n28) );
  AOI22_X1 OutputReg_U47 ( .A1(OutputReg_n69), .A2(Output[26]), .B1(
        OutputReg_n2), .B2(OutputRegIn[26]), .ZN(OutputReg_n29) );
  AOI22_X1 OutputReg_U46 ( .A1(OutputReg_n69), .A2(Output[27]), .B1(
        OutputReg_n3), .B2(OutputRegIn[27]), .ZN(OutputReg_n30) );
  AOI22_X1 OutputReg_U45 ( .A1(OutputReg_n69), .A2(Output[28]), .B1(
        OutputReg_n67), .B2(OutputRegIn[28]), .ZN(OutputReg_n31) );
  AOI22_X1 OutputReg_U44 ( .A1(OutputReg_n69), .A2(Output[29]), .B1(
        OutputReg_n67), .B2(OutputRegIn[29]), .ZN(OutputReg_n32) );
  AOI22_X1 OutputReg_U43 ( .A1(OutputReg_n69), .A2(Output[30]), .B1(
        OutputReg_n67), .B2(OutputRegIn[30]), .ZN(OutputReg_n33) );
  AOI22_X1 OutputReg_U42 ( .A1(OutputReg_n69), .A2(Output[31]), .B1(
        OutputReg_n67), .B2(OutputRegIn[31]), .ZN(OutputReg_n34) );
  AOI22_X1 OutputReg_U41 ( .A1(OutputReg_n69), .A2(Output[32]), .B1(
        OutputReg_n67), .B2(OutputRegIn[32]), .ZN(OutputReg_n35) );
  AOI22_X1 OutputReg_U40 ( .A1(OutputReg_n69), .A2(Output[33]), .B1(
        OutputReg_n67), .B2(OutputRegIn[33]), .ZN(OutputReg_n36) );
  AOI22_X1 OutputReg_U39 ( .A1(OutputReg_n71), .A2(Output[34]), .B1(
        OutputReg_n67), .B2(OutputRegIn[34]), .ZN(OutputReg_n37) );
  AOI22_X1 OutputReg_U38 ( .A1(OutputReg_n71), .A2(Output[35]), .B1(
        OutputReg_n67), .B2(OutputRegIn[35]), .ZN(OutputReg_n38) );
  AOI22_X1 OutputReg_U37 ( .A1(OutputReg_n71), .A2(Output[36]), .B1(
        OutputReg_n67), .B2(OutputRegIn[36]), .ZN(OutputReg_n39) );
  AOI22_X1 OutputReg_U36 ( .A1(OutputReg_n71), .A2(Output[37]), .B1(
        OutputReg_n67), .B2(OutputRegIn[37]), .ZN(OutputReg_n40) );
  AOI22_X1 OutputReg_U35 ( .A1(OutputReg_n71), .A2(Output[38]), .B1(
        OutputReg_n67), .B2(OutputRegIn[38]), .ZN(OutputReg_n41) );
  AOI22_X1 OutputReg_U34 ( .A1(OutputReg_n71), .A2(Output[39]), .B1(
        OutputReg_n67), .B2(OutputRegIn[39]), .ZN(OutputReg_n42) );
  AOI22_X1 OutputReg_U33 ( .A1(OutputReg_n71), .A2(Output[40]), .B1(
        OutputReg_n3), .B2(OutputRegIn[40]), .ZN(OutputReg_n43) );
  AOI22_X1 OutputReg_U32 ( .A1(OutputReg_n68), .A2(Output[41]), .B1(
        OutputReg_n3), .B2(OutputRegIn[41]), .ZN(OutputReg_n44) );
  AOI22_X1 OutputReg_U31 ( .A1(OutputReg_n68), .A2(Output[42]), .B1(
        OutputReg_n3), .B2(OutputRegIn[42]), .ZN(OutputReg_n45) );
  AOI22_X1 OutputReg_U30 ( .A1(OutputReg_n68), .A2(Output[43]), .B1(
        OutputReg_n3), .B2(OutputRegIn[43]), .ZN(OutputReg_n46) );
  AOI22_X1 OutputReg_U29 ( .A1(OutputReg_n68), .A2(Output[44]), .B1(
        OutputReg_n3), .B2(OutputRegIn[44]), .ZN(OutputReg_n47) );
  AOI22_X1 OutputReg_U28 ( .A1(OutputReg_n68), .A2(Output[45]), .B1(
        OutputReg_n3), .B2(OutputRegIn[45]), .ZN(OutputReg_n48) );
  AOI22_X1 OutputReg_U27 ( .A1(OutputReg_n68), .A2(Output[46]), .B1(
        OutputReg_n3), .B2(OutputRegIn[46]), .ZN(OutputReg_n49) );
  AOI22_X1 OutputReg_U26 ( .A1(OutputReg_n68), .A2(Output[47]), .B1(
        OutputReg_n3), .B2(OutputRegIn[47]), .ZN(OutputReg_n50) );
  AOI22_X1 OutputReg_U25 ( .A1(OutputReg_n68), .A2(Output[48]), .B1(
        OutputReg_n3), .B2(OutputRegIn[48]), .ZN(OutputReg_n51) );
  AOI22_X1 OutputReg_U24 ( .A1(OutputReg_n68), .A2(Output[49]), .B1(
        OutputReg_n3), .B2(OutputRegIn[49]), .ZN(OutputReg_n52) );
  AOI22_X1 OutputReg_U23 ( .A1(OutputReg_n68), .A2(Output[50]), .B1(
        OutputReg_n3), .B2(OutputRegIn[50]), .ZN(OutputReg_n53) );
  AOI22_X1 OutputReg_U22 ( .A1(OutputReg_n68), .A2(Output[51]), .B1(
        OutputReg_n3), .B2(OutputRegIn[51]), .ZN(OutputReg_n54) );
  AOI22_X1 OutputReg_U21 ( .A1(OutputReg_n68), .A2(Output[52]), .B1(
        OutputReg_n2), .B2(OutputRegIn[52]), .ZN(OutputReg_n55) );
  AOI22_X1 OutputReg_U20 ( .A1(OutputReg_n68), .A2(Output[53]), .B1(
        OutputReg_n2), .B2(OutputRegIn[53]), .ZN(OutputReg_n56) );
  AOI22_X1 OutputReg_U19 ( .A1(OutputReg_n68), .A2(Output[54]), .B1(
        OutputReg_n2), .B2(OutputRegIn[54]), .ZN(OutputReg_n57) );
  AOI22_X1 OutputReg_U18 ( .A1(OutputReg_n68), .A2(Output[55]), .B1(
        OutputReg_n2), .B2(OutputRegIn[55]), .ZN(OutputReg_n58) );
  AOI22_X1 OutputReg_U17 ( .A1(OutputReg_n68), .A2(Output[56]), .B1(
        OutputReg_n2), .B2(OutputRegIn[56]), .ZN(OutputReg_n59) );
  AOI22_X1 OutputReg_U16 ( .A1(OutputReg_n68), .A2(Output[57]), .B1(
        OutputReg_n2), .B2(OutputRegIn[57]), .ZN(OutputReg_n60) );
  AOI22_X1 OutputReg_U15 ( .A1(OutputReg_n68), .A2(Output[58]), .B1(
        OutputReg_n2), .B2(OutputRegIn[58]), .ZN(OutputReg_n61) );
  AOI22_X1 OutputReg_U14 ( .A1(OutputReg_n68), .A2(Output[59]), .B1(
        OutputReg_n2), .B2(OutputRegIn[59]), .ZN(OutputReg_n62) );
  AOI22_X1 OutputReg_U13 ( .A1(OutputReg_n68), .A2(Output[60]), .B1(
        OutputReg_n2), .B2(OutputRegIn[60]), .ZN(OutputReg_n63) );
  AOI22_X1 OutputReg_U12 ( .A1(OutputReg_n68), .A2(Output[61]), .B1(
        OutputReg_n2), .B2(OutputRegIn[61]), .ZN(OutputReg_n64) );
  AOI22_X1 OutputReg_U11 ( .A1(OutputReg_n68), .A2(Output[62]), .B1(
        OutputReg_n2), .B2(OutputRegIn[62]), .ZN(OutputReg_n65) );
  AOI22_X1 OutputReg_U10 ( .A1(OutputReg_n68), .A2(Output[63]), .B1(
        OutputReg_n2), .B2(OutputRegIn[63]), .ZN(OutputReg_n66) );
  NOR2_X1 OutputReg_U9 ( .A1(done), .A2(rst), .ZN(OutputReg_n71) );
  BUF_X1 OutputReg_U8 ( .A(OutputReg_n71), .Z(OutputReg_n69) );
  BUF_X2 OutputReg_U7 ( .A(OutputReg_n71), .Z(OutputReg_n68) );
  NOR2_X1 OutputReg_U6 ( .A1(rst), .A2(OutputReg_n68), .ZN(OutputReg_n70) );
  BUF_X1 OutputReg_U5 ( .A(OutputReg_n70), .Z(OutputReg_n3) );
  BUF_X1 OutputReg_U4 ( .A(OutputReg_n70), .Z(OutputReg_n2) );
  BUF_X1 OutputReg_U3 ( .A(OutputReg_n70), .Z(OutputReg_n67) );
  DFF_X1 OutputReg_Q_reg_0_ ( .D(OutputReg_n1), .CK(clk), .Q(), .QN(Output[0])
         );
  DFF_X1 OutputReg_Q_reg_1_ ( .D(OutputReg_n4), .CK(clk), .Q(), .QN(Output[1])
         );
  DFF_X1 OutputReg_Q_reg_2_ ( .D(OutputReg_n5), .CK(clk), .Q(), .QN(Output[2])
         );
  DFF_X1 OutputReg_Q_reg_3_ ( .D(OutputReg_n6), .CK(clk), .Q(), .QN(Output[3])
         );
  DFF_X1 OutputReg_Q_reg_4_ ( .D(OutputReg_n7), .CK(clk), .Q(), .QN(Output[4])
         );
  DFF_X1 OutputReg_Q_reg_5_ ( .D(OutputReg_n8), .CK(clk), .Q(), .QN(Output[5])
         );
  DFF_X1 OutputReg_Q_reg_6_ ( .D(OutputReg_n9), .CK(clk), .Q(), .QN(Output[6])
         );
  DFF_X1 OutputReg_Q_reg_7_ ( .D(OutputReg_n10), .CK(clk), .Q(), .QN(Output[7]) );
  DFF_X1 OutputReg_Q_reg_8_ ( .D(OutputReg_n11), .CK(clk), .Q(), .QN(Output[8]) );
  DFF_X1 OutputReg_Q_reg_9_ ( .D(OutputReg_n12), .CK(clk), .Q(), .QN(Output[9]) );
  DFF_X1 OutputReg_Q_reg_10_ ( .D(OutputReg_n13), .CK(clk), .Q(), .QN(
        Output[10]) );
  DFF_X1 OutputReg_Q_reg_11_ ( .D(OutputReg_n14), .CK(clk), .Q(), .QN(
        Output[11]) );
  DFF_X1 OutputReg_Q_reg_12_ ( .D(OutputReg_n15), .CK(clk), .Q(), .QN(
        Output[12]) );
  DFF_X1 OutputReg_Q_reg_13_ ( .D(OutputReg_n16), .CK(clk), .Q(), .QN(
        Output[13]) );
  DFF_X1 OutputReg_Q_reg_14_ ( .D(OutputReg_n17), .CK(clk), .Q(), .QN(
        Output[14]) );
  DFF_X1 OutputReg_Q_reg_15_ ( .D(OutputReg_n18), .CK(clk), .Q(), .QN(
        Output[15]) );
  DFF_X1 OutputReg_Q_reg_16_ ( .D(OutputReg_n19), .CK(clk), .Q(), .QN(
        Output[16]) );
  DFF_X1 OutputReg_Q_reg_17_ ( .D(OutputReg_n20), .CK(clk), .Q(), .QN(
        Output[17]) );
  DFF_X1 OutputReg_Q_reg_18_ ( .D(OutputReg_n21), .CK(clk), .Q(), .QN(
        Output[18]) );
  DFF_X1 OutputReg_Q_reg_19_ ( .D(OutputReg_n22), .CK(clk), .Q(), .QN(
        Output[19]) );
  DFF_X1 OutputReg_Q_reg_20_ ( .D(OutputReg_n23), .CK(clk), .Q(), .QN(
        Output[20]) );
  DFF_X1 OutputReg_Q_reg_21_ ( .D(OutputReg_n24), .CK(clk), .Q(), .QN(
        Output[21]) );
  DFF_X1 OutputReg_Q_reg_22_ ( .D(OutputReg_n25), .CK(clk), .Q(), .QN(
        Output[22]) );
  DFF_X1 OutputReg_Q_reg_23_ ( .D(OutputReg_n26), .CK(clk), .Q(), .QN(
        Output[23]) );
  DFF_X1 OutputReg_Q_reg_24_ ( .D(OutputReg_n27), .CK(clk), .Q(), .QN(
        Output[24]) );
  DFF_X1 OutputReg_Q_reg_25_ ( .D(OutputReg_n28), .CK(clk), .Q(), .QN(
        Output[25]) );
  DFF_X1 OutputReg_Q_reg_26_ ( .D(OutputReg_n29), .CK(clk), .Q(), .QN(
        Output[26]) );
  DFF_X1 OutputReg_Q_reg_27_ ( .D(OutputReg_n30), .CK(clk), .Q(), .QN(
        Output[27]) );
  DFF_X1 OutputReg_Q_reg_28_ ( .D(OutputReg_n31), .CK(clk), .Q(), .QN(
        Output[28]) );
  DFF_X1 OutputReg_Q_reg_29_ ( .D(OutputReg_n32), .CK(clk), .Q(), .QN(
        Output[29]) );
  DFF_X1 OutputReg_Q_reg_30_ ( .D(OutputReg_n33), .CK(clk), .Q(), .QN(
        Output[30]) );
  DFF_X1 OutputReg_Q_reg_31_ ( .D(OutputReg_n34), .CK(clk), .Q(), .QN(
        Output[31]) );
  DFF_X1 OutputReg_Q_reg_32_ ( .D(OutputReg_n35), .CK(clk), .Q(), .QN(
        Output[32]) );
  DFF_X1 OutputReg_Q_reg_33_ ( .D(OutputReg_n36), .CK(clk), .Q(), .QN(
        Output[33]) );
  DFF_X1 OutputReg_Q_reg_34_ ( .D(OutputReg_n37), .CK(clk), .Q(), .QN(
        Output[34]) );
  DFF_X1 OutputReg_Q_reg_35_ ( .D(OutputReg_n38), .CK(clk), .Q(), .QN(
        Output[35]) );
  DFF_X1 OutputReg_Q_reg_36_ ( .D(OutputReg_n39), .CK(clk), .Q(), .QN(
        Output[36]) );
  DFF_X1 OutputReg_Q_reg_37_ ( .D(OutputReg_n40), .CK(clk), .Q(), .QN(
        Output[37]) );
  DFF_X1 OutputReg_Q_reg_38_ ( .D(OutputReg_n41), .CK(clk), .Q(), .QN(
        Output[38]) );
  DFF_X1 OutputReg_Q_reg_39_ ( .D(OutputReg_n42), .CK(clk), .Q(), .QN(
        Output[39]) );
  DFF_X1 OutputReg_Q_reg_40_ ( .D(OutputReg_n43), .CK(clk), .Q(), .QN(
        Output[40]) );
  DFF_X1 OutputReg_Q_reg_41_ ( .D(OutputReg_n44), .CK(clk), .Q(), .QN(
        Output[41]) );
  DFF_X1 OutputReg_Q_reg_42_ ( .D(OutputReg_n45), .CK(clk), .Q(), .QN(
        Output[42]) );
  DFF_X1 OutputReg_Q_reg_43_ ( .D(OutputReg_n46), .CK(clk), .Q(), .QN(
        Output[43]) );
  DFF_X1 OutputReg_Q_reg_44_ ( .D(OutputReg_n47), .CK(clk), .Q(), .QN(
        Output[44]) );
  DFF_X1 OutputReg_Q_reg_45_ ( .D(OutputReg_n48), .CK(clk), .Q(), .QN(
        Output[45]) );
  DFF_X1 OutputReg_Q_reg_46_ ( .D(OutputReg_n49), .CK(clk), .Q(), .QN(
        Output[46]) );
  DFF_X1 OutputReg_Q_reg_47_ ( .D(OutputReg_n50), .CK(clk), .Q(), .QN(
        Output[47]) );
  DFF_X1 OutputReg_Q_reg_48_ ( .D(OutputReg_n51), .CK(clk), .Q(), .QN(
        Output[48]) );
  DFF_X1 OutputReg_Q_reg_49_ ( .D(OutputReg_n52), .CK(clk), .Q(), .QN(
        Output[49]) );
  DFF_X1 OutputReg_Q_reg_50_ ( .D(OutputReg_n53), .CK(clk), .Q(), .QN(
        Output[50]) );
  DFF_X1 OutputReg_Q_reg_51_ ( .D(OutputReg_n54), .CK(clk), .Q(), .QN(
        Output[51]) );
  DFF_X1 OutputReg_Q_reg_52_ ( .D(OutputReg_n55), .CK(clk), .Q(), .QN(
        Output[52]) );
  DFF_X1 OutputReg_Q_reg_53_ ( .D(OutputReg_n56), .CK(clk), .Q(), .QN(
        Output[53]) );
  DFF_X1 OutputReg_Q_reg_54_ ( .D(OutputReg_n57), .CK(clk), .Q(), .QN(
        Output[54]) );
  DFF_X1 OutputReg_Q_reg_55_ ( .D(OutputReg_n58), .CK(clk), .Q(), .QN(
        Output[55]) );
  DFF_X1 OutputReg_Q_reg_56_ ( .D(OutputReg_n59), .CK(clk), .Q(), .QN(
        Output[56]) );
  DFF_X1 OutputReg_Q_reg_57_ ( .D(OutputReg_n60), .CK(clk), .Q(), .QN(
        Output[57]) );
  DFF_X1 OutputReg_Q_reg_58_ ( .D(OutputReg_n61), .CK(clk), .Q(), .QN(
        Output[58]) );
  DFF_X1 OutputReg_Q_reg_59_ ( .D(OutputReg_n62), .CK(clk), .Q(), .QN(
        Output[59]) );
  DFF_X1 OutputReg_Q_reg_60_ ( .D(OutputReg_n63), .CK(clk), .Q(), .QN(
        Output[60]) );
  DFF_X1 OutputReg_Q_reg_61_ ( .D(OutputReg_n64), .CK(clk), .Q(), .QN(
        Output[61]) );
  DFF_X1 OutputReg_Q_reg_62_ ( .D(OutputReg_n65), .CK(clk), .Q(), .QN(
        Output[62]) );
  DFF_X1 OutputReg_Q_reg_63_ ( .D(OutputReg_n66), .CK(clk), .Q(), .QN(
        Output[63]) );
endmodule

